
module c5315_synth ( N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, 
        N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, 
        N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, 
        N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, 
        N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, 
        N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, 
        N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, 
        N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, 
        N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, 
        N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, 
        N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, 
        N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, 
        N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, 
        N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, 
        N610, N613, N616, N619, N625, N631, N709, N816, N1066, N1137, N1138, 
        N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, 
        N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, 
        N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, 
        N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, 
        N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, 
        N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, 
        N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, 
        N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, 
        N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, 
        N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, 
        N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, 
        N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128 );
  input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37,
         N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79,
         N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106,
         N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136,
         N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164,
         N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197,
         N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234,
         N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273,
         N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315,
         N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358,
         N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422,
         N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545,
         N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583,
         N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610,
         N613, N616, N619, N625, N631;
  output N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060,
         N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357,
         N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737,
         N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716,
         N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449,
         N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476,
         N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520,
         N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607,
         N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706,
         N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754,
         N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123,
         N8124, N8127, N8128;
  wire   N1042, N1043, N1067, N1080, N1092, N1104, N1146, N1148, N1149, N1150,
         N1151, N1156, N1157, N1161, N1173, N1185, N1197, N1209, N1213, N1216,
         N1219, N1223, N1235, N1247, N1259, N1271, N1280, N1292, N1303, N1315,
         N1327, N1339, N1351, N1363, N1375, N1378, N1381, N1384, N1387, N1390,
         N1393, N1396, N1415, N1418, N1421, N1424, N1427, N1430, N1433, N1436,
         N1455, N1462, N1469, N1475, N1479, N1482, N1492, N1495, N1498, N1501,
         N1504, N1507, N1510, N1513, N1516, N1519, N1522, N1525, N1542, N1545,
         N1548, N1551, N1554, N1557, N1560, N1563, N1566, N1573, N1580, N1583,
         N1588, N1594, N1597, N1600, N1603, N1606, N1609, N1612, N1615, N1618,
         N1621, N1624, N1627, N1630, N1633, N1636, N1639, N1642, N1645, N1648,
         N1651, N1654, N1657, N1660, N1663, N1675, N1685, N1697, N1709, N1721,
         N1727, N1731, N1743, N1755, N1758, N1761, N1769, N1777, N1785, N1793,
         N1800, N1807, N1814, N1821, N1824, N1827, N1830, N1833, N1836, N1839,
         N1842, N1845, N1848, N1851, N1854, N1857, N1860, N1863, N1866, N1869,
         N1872, N1875, N1878, N1881, N1884, N1887, N1890, N1893, N1896, N1899,
         N1902, N1905, N1908, N1911, N1914, N1917, N1920, N1923, N1926, N1929,
         N1932, N1935, N1938, N1941, N1944, N1947, N1950, N1953, N1956, N1959,
         N1962, N1965, N1968, N2349, N2350, N2585, N2586, N2587, N2588, N2589,
         N2591, N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599, N2600,
         N2601, N2602, N2603, N2604, N2605, N2606, N2607, N2608, N2609, N2610,
         N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619, N2620,
         N2621, N2622, N2624, N2625, N2626, N2627, N2628, N2629, N2630, N2631,
         N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641,
         N2642, N2643, N2644, N2645, N2646, N2647, N2653, N2664, N2675, N2681,
         N2692, N2703, N2704, N2709, N2710, N2711, N2712, N2713, N2714, N2715,
         N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2728, N2739, N2750,
         N2756, N2767, N2778, N2779, N2790, N2801, N2812, N2823, N2824, N2825,
         N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835,
         N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845,
         N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855,
         N2861, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875,
         N2876, N2877, N2882, N2891, N2901, N2902, N2903, N2904, N2905, N2906,
         N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916,
         N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926,
         N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936,
         N2937, N2938, N2939, N2940, N2941, N2942, N2948, N2954, N2955, N2956,
         N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2969, N2970,
         N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979, N2980,
         N2981, N2982, N2983, N2984, N2985, N2986, N2987, N2988, N2989, N2990,
         N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000,
         N3003, N3006, N3007, N3010, N3013, N3014, N3015, N3016, N3017, N3018,
         N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028,
         N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3038, N3041, N3052,
         N3063, N3068, N3071, N3072, N3073, N3074, N3075, N3086, N3097, N3108,
         N3119, N3130, N3141, N3142, N3143, N3144, N3145, N3146, N3147, N3158,
         N3169, N3180, N3191, N3194, N3195, N3196, N3197, N3198, N3199, N3200,
         N3203, N3401, N3402, N3403, N3404, N3405, N3406, N3407, N3408, N3409,
         N3410, N3411, N3412, N3413, N3414, N3415, N3416, N3444, N3445, N3446,
         N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456,
         N3459, N3460, N3461, N3462, N3463, N3464, N3465, N3466, N3481, N3482,
         N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492,
         N3493, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510,
         N3511, N3512, N3513, N3514, N3515, N3558, N3559, N3560, N3561, N3562,
         N3563, N3605, N3606, N3607, N3608, N3609, N3610, N3614, N3615, N3616,
         N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, N3625, N3626,
         N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636,
         N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, N3645, N3646,
         N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656,
         N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3665, N3666,
         N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676,
         N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686,
         N3687, N3688, N3689, N3691, N3700, N3701, N3702, N3703, N3704, N3705,
         N3708, N3709, N3710, N3711, N3712, N3713, N3715, N3716, N3717, N3718,
         N3719, N3720, N3721, N3722, N3723, N3724, N3725, N3726, N3727, N3728,
         N3729, N3730, N3731, N3732, N3738, N3739, N3740, N3741, N3742, N3743,
         N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753,
         N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763,
         N3764, N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3775, N3779,
         N3780, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3789,
         N3793, N3797, N3800, N3801, N3802, N3803, N3804, N3805, N3806, N3807,
         N3808, N3809, N3810, N3813, N3816, N3819, N3822, N3823, N3824, N3827,
         N3828, N3829, N3830, N3831, N3834, N3835, N3836, N3837, N3838, N3839,
         N3840, N3841, N3842, N3849, N3855, N3861, N3867, N3873, N3881, N3887,
         N3893, N3908, N3909, N3911, N3914, N3915, N3916, N3917, N3918, N3919,
         N3920, N3921, N3927, N3933, N3942, N3948, N3956, N3962, N3968, N3975,
         N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, N3987,
         N3988, N3989, N3990, N3991, N3998, N4008, N4011, N4021, N4024, N4027,
         N4031, N4032, N4033, N4034, N4035, N4036, N4037, N4038, N4039, N4040,
         N4041, N4042, N4067, N4080, N4088, N4091, N4094, N4097, N4100, N4103,
         N4106, N4109, N4144, N4147, N4150, N4153, N4156, N4159, N4183, N4184,
         N4185, N4186, N4188, N4191, N4196, N4197, N4198, N4199, N4200, N4203,
         N4206, N4209, N4212, N4215, N4219, N4223, N4224, N4225, N4228, N4231,
         N4234, N4237, N4240, N4243, N4246, N4249, N4252, N4255, N4258, N4263,
         N4264, N4267, N4268, N4269, N4270, N4271, N4273, N4274, N4276, N4277,
         N4280, N4284, N4290, N4297, N4298, N4301, N4305, N4310, N4316, N4320,
         N4325, N4331, N4332, N4336, N4342, N4349, N4357, N4364, N4375, N4379,
         N4385, N4392, N4396, N4400, N4405, N4412, N4418, N4425, N4436, N4440,
         N4445, N4451, N4456, N4462, N4469, N4477, N4512, N4515, N4516, N4521,
         N4523, N4524, N4532, N4547, N4548, N4551, N4554, N4557, N4560, N4563,
         N4566, N4569, N4572, N4575, N4578, N4581, N4584, N4587, N4590, N4593,
         N4596, N4599, N4602, N4605, N4608, N4611, N4614, N4617, N4621, N4624,
         N4627, N4630, N4633, N4637, N4640, N4643, N4646, N4649, N4652, N4655,
         N4658, N4662, N4665, N4668, N4671, N4674, N4677, N4680, N4683, N4686,
         N4689, N4692, N4695, N4698, N4701, N4702, N4720, N4721, N4724, N4725,
         N4726, N4727, N4728, N4729, N4730, N4731, N4732, N4733, N4734, N4735,
         N4736, N4741, N4855, N4856, N4908, N4909, N4939, N4942, N4947, N4953,
         N4954, N4955, N4956, N4957, N4958, N4959, N4960, N4961, N4965, N4966,
         N4967, N4968, N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979,
         N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N5049, N5052,
         N5053, N5054, N5055, N5056, N5057, N5058, N5059, N5060, N5061, N5062,
         N5063, N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073,
         N5074, N5075, N5076, N5077, N5078, N5079, N5080, N5081, N5082, N5083,
         N5084, N5085, N5086, N5087, N5088, N5089, N5090, N5091, N5092, N5093,
         N5094, N5095, N5096, N5097, N5098, N5099, N5100, N5101, N5102, N5103,
         N5104, N5105, N5106, N5107, N5108, N5109, N5110, N5111, N5112, N5113,
         N5114, N5115, N5116, N5117, N5118, N5119, N5120, N5121, N5122, N5123,
         N5124, N5125, N5126, N5127, N5128, N5129, N5130, N5131, N5132, N5133,
         N5135, N5136, N5137, N5138, N5139, N5140, N5141, N5142, N5143, N5144,
         N5145, N5146, N5147, N5148, N5150, N5153, N5154, N5155, N5156, N5157,
         N5160, N5161, N5162, N5163, N5164, N5165, N5166, N5169, N5172, N5173,
         N5176, N5177, N5180, N5183, N5186, N5189, N5192, N5195, N5198, N5199,
         N5202, N5205, N5208, N5211, N5214, N5217, N5220, N5223, N5224, N5225,
         N5226, N5227, N5228, N5229, N5230, N5232, N5233, N5234, N5235, N5236,
         N5239, N5241, N5242, N5243, N5244, N5245, N5246, N5247, N5248, N5249,
         N5250, N5252, N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260,
         N5261, N5262, N5263, N5264, N5274, N5275, N5282, N5283, N5284, N5298,
         N5299, N5300, N5303, N5304, N5305, N5306, N5307, N5308, N5309, N5310,
         N5311, N5312, N5315, N5319, N5324, N5328, N5331, N5332, N5346, N5363,
         N5364, N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5374, N5377,
         N5382, N5385, N5389, N5396, N5407, N5418, N5424, N5431, N5441, N5452,
         N5462, N5469, N5470, N5477, N5488, N5498, N5506, N5520, N5536, N5549,
         N5555, N5562, N5573, N5579, N5595, N5606, N5616, N5617, N5618, N5619,
         N5620, N5621, N5622, N5624, N5634, N5655, N5671, N5684, N5690, N5691,
         N5692, N5696, N5700, N5703, N5707, N5711, N5726, N5727, N5728, N5730,
         N5731, N5732, N5733, N5734, N5735, N5736, N5739, N5742, N5745, N5755,
         N5756, N5954, N5955, N5956, N6005, N6006, N6023, N6024, N6025, N6028,
         N6031, N6034, N6037, N6040, N6044, N6045, N6048, N6051, N6054, N6065,
         N6066, N6067, N6068, N6069, N6071, N6072, N6073, N6074, N6075, N6076,
         N6077, N6078, N6079, N6080, N6083, N6084, N6085, N6086, N6087, N6088,
         N6089, N6090, N6091, N6094, N6095, N6096, N6097, N6098, N6099, N6100,
         N6101, N6102, N6103, N6104, N6105, N6106, N6107, N6108, N6111, N6112,
         N6113, N6114, N6115, N6116, N6117, N6120, N6121, N6122, N6123, N6124,
         N6125, N6126, N6127, N6128, N6129, N6130, N6131, N6132, N6133, N6134,
         N6135, N6136, N6137, N6138, N6139, N6140, N6143, N6144, N6145, N6146,
         N6147, N6148, N6149, N6152, N6153, N6154, N6155, N6156, N6157, N6158,
         N6159, N6160, N6161, N6162, N6163, N6164, N6168, N6171, N6172, N6173,
         N6174, N6175, N6178, N6179, N6180, N6181, N6182, N6183, N6184, N6185,
         N6186, N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6197,
         N6200, N6203, N6206, N6209, N6212, N6215, N6218, N6221, N6234, N6235,
         N6238, N6241, N6244, N6247, N6250, N6253, N6256, N6259, N6262, N6265,
         N6268, N6271, N6274, N6277, N6280, N6283, N6286, N6289, N6292, N6295,
         N6298, N6301, N6304, N6307, N6310, N6313, N6316, N6319, N6322, N6325,
         N6328, N6331, N6335, N6338, N6341, N6344, N6347, N6350, N6353, N6356,
         N6359, N6364, N6367, N6370, N6373, N6374, N6375, N6376, N6377, N6378,
         N6382, N6386, N6388, N6392, N6397, N6411, N6415, N6419, N6427, N6434,
         N6437, N6441, N6445, N6448, N6449, N6466, N6469, N6470, N6471, N6472,
         N6473, N6474, N6475, N6476, N6477, N6478, N6482, N6486, N6490, N6494,
         N6500, N6504, N6508, N6512, N6516, N6526, N6536, N6539, N6553, N6556,
         N6566, N6569, N6572, N6575, N6580, N6584, N6587, N6592, N6599, N6606,
         N6609, N6619, N6622, N6630, N6631, N6632, N6633, N6634, N6637, N6640,
         N6650, N6651, N6653, N6655, N6657, N6659, N6660, N6661, N6662, N6663,
         N6664, N6666, N6668, N6670, N6672, N6675, N6680, N6681, N6682, N6683,
         N6689, N6690, N6691, N6692, N6693, N6695, N6698, N6699, N6700, N6703,
         N6708, N6709, N6710, N6711, N6712, N6713, N6714, N6715, N6718, N6719,
         N6720, N6721, N6722, N6724, N6739, N6740, N6741, N6744, N6745, N6746,
         N6751, N6752, N6753, N6754, N6755, N6760, N6761, N6762, N6772, N6773,
         N6776, N6777, N6782, N6783, N6784, N6785, N6790, N6791, N6792, N6795,
         N6801, N6802, N6803, N6804, N6805, N6806, N6807, N6808, N6809, N6810,
         N6811, N6812, N6813, N6814, N6815, N6816, N6817, N6823, N6824, N6825,
         N6826, N6827, N6828, N6829, N6830, N6831, N6834, N6835, N6836, N6837,
         N6838, N6839, N6840, N6841, N6842, N6843, N6844, N6850, N6851, N6852,
         N6853, N6854, N6855, N6856, N6857, N6860, N6861, N6862, N6863, N6866,
         N6872, N6873, N6874, N6875, N6876, N6879, N6880, N6881, N6884, N6885,
         N6888, N6889, N6890, N6891, N6894, N6895, N6896, N6897, N6900, N6901,
         N6904, N6905, N6908, N6909, N6912, N6913, N6914, N6915, N6916, N6919,
         N6922, N6923, N6930, N6932, N6935, N6936, N6937, N6938, N6939, N6940,
         N6946, N6947, N6948, N6949, N6953, N6954, N6955, N6956, N6957, N6958,
         N6964, N6965, N6966, N6967, N6973, N6974, N6975, N6976, N6977, N6978,
         N6979, N6987, N6990, N6999, N7002, N7003, N7006, N7011, N7012, N7013,
         N7016, N7018, N7019, N7020, N7021, N7022, N7023, N7028, N7031, N7034,
         N7037, N7040, N7041, N7044, N7045, N7046, N7047, N7048, N7049, N7054,
         N7057, N7060, N7064, N7065, N7072, N7073, N7074, N7075, N7076, N7079,
         N7080, N7083, N7084, N7085, N7086, N7087, N7088, N7089, N7090, N7093,
         N7094, N7097, N7101, N7105, N7110, N7114, N7115, N7116, N7125, N7126,
         N7127, N7130, N7131, N7139, N7140, N7141, N7146, N7147, N7149, N7150,
         N7151, N7152, N7153, N7158, N7159, N7160, N7166, N7167, N7168, N7169,
         N7170, N7171, N7172, N7173, N7174, N7175, N7176, N7177, N7178, N7179,
         N7180, N7181, N7182, N7183, N7184, N7185, N7186, N7187, N7188, N7189,
         N7190, N7196, N7197, N7198, N7204, N7205, N7206, N7207, N7208, N7209,
         N7212, N7215, N7216, N7217, N7218, N7219, N7222, N7225, N7228, N7229,
         N7236, N7239, N7242, N7245, N7250, N7257, N7260, N7263, N7268, N7269,
         N7270, N7276, N7282, N7288, N7294, N7300, N7301, N7304, N7310, N7320,
         N7321, N7328, N7338, N7339, N7340, N7341, N7342, N7349, N7357, N7364,
         N7394, N7397, N7402, N7405, N7406, N7407, N7408, N7409, N7412, N7415,
         N7416, N7417, N7418, N7419, N7420, N7421, N7424, N7425, N7426, N7427,
         N7428, N7429, N7430, N7431, N7433, N7434, N7435, N7436, N7437, N7438,
         N7439, N7440, N7441, N7442, N7443, N7444, N7445, N7446, N7447, N7448,
         N7450, N7451, N7452, N7453, N7454, N7455, N7456, N7457, N7458, N7459,
         N7460, N7461, N7462, N7463, N7464, N7468, N7479, N7481, N7482, N7483,
         N7484, N7485, N7486, N7487, N7488, N7489, N7492, N7493, N7498, N7499,
         N7500, N7505, N7507, N7508, N7509, N7510, N7512, N7513, N7514, N7525,
         N7526, N7527, N7528, N7529, N7530, N7531, N7537, N7543, N7549, N7555,
         N7561, N7567, N7573, N7579, N7582, N7585, N7586, N7587, N7588, N7589,
         N7592, N7595, N7598, N7599, N7624, N7625, N7631, N7636, N7657, N7658,
         N7665, N7666, N7667, N7668, N7669, N7670, N7671, N7672, N7673, N7674,
         N7675, N7676, N7677, N7678, N7679, N7680, N7681, N7682, N7683, N7684,
         N7685, N7686, N7687, N7688, N7689, N7690, N7691, N7692, N7693, N7694,
         N7695, N7696, N7697, N7708, N7709, N7710, N7711, N7712, N7715, N7718,
         N7719, N7720, N7721, N7722, N7723, N7724, N7727, N7728, N7729, N7730,
         N7731, N7732, N7733, N7734, N7743, N7744, N7749, N7750, N7751, N7762,
         N7765, N7768, N7769, N7770, N7771, N7772, N7775, N7778, N7781, N7782,
         N7787, N7788, N7795, N7796, N7797, N7798, N7799, N7800, N7803, N7806,
         N7807, N7808, N7809, N7810, N7811, N7812, N7815, N7816, N7821, N7822,
         N7823, N7826, N7829, N7832, N7833, N7834, N7835, N7836, N7839, N7842,
         N7845, N7846, N7851, N7852, N7859, N7860, N7861, N7862, N7863, N7864,
         N7867, N7870, N7871, N7872, N7873, N7874, N7875, N7876, N7879, N7880,
         N7885, N7886, N7887, N7890, N7893, N7896, N7897, N7898, N7899, N7900,
         N7903, N7906, N7909, N7910, N7917, N7918, N7923, N7924, N7925, N7926,
         N7927, N7928, N7929, N7930, N7931, N7932, N7935, N7938, N7939, N7940,
         N7943, N7944, N7945, N7946, N7951, N7954, N7957, N7960, N7963, N7966,
         N7967, N7968, N7969, N7970, N7973, N7974, N7984, N7985, N7987, N7988,
         N7989, N7990, N7991, N7992, N7993, N7994, N7995, N7996, N7997, N7998,
         N8001, N8004, N8009, N8013, N8017, N8020, N8021, N8022, N8023, N8025,
         N8026, N8027, N8031, N8032, N8033, N8034, N8035, N8036, N8037, N8038,
         N8039, N8040, N8041, N8042, N8043, N8044, N8045, N8048, N8055, N8056,
         N8057, N8058, N8059, N8060, N8061, N8064, N8071, N8072, N8073, N8074,
         N8077, N8078, N8079, N8082, N8089, N8090, N8091, N8092, N8093, N8096,
         N8099, N8102, N8113, N8114, N8115, N8116, N8117, N8118, N8119, N8120,
         N8121, N8122, N8125, N8126, N1156_1, N1156_2, N2585_1, N2586_1,
         N2587_1, N2588_1, N2589_1, N2591_1, N2592_1, N2593_1, N2594_1,
         N2595_1, N2596_1, N2597_1, N2598_1, N2599_1, N2600_1, N2601_1,
         N2602_1, N2603_1, N2604_1, N2605_1, N2606_1, N2607_1, N2608_1,
         N2609_1, N2610_1, N2611_1, N2612_1, N2613_1, N2614_1, N2615_1,
         N2616_1, N2617_1, N2618_1, N2619_1, N2620_1, N2621_1, N2622_1,
         N2624_1, N2626_1, N2703_1, N2778_1, N2831_1, N2832_1, N2833_1,
         N2834_1, N2847_1, N2848_1, N2849_1, N2850_1, N2908_1, N2909_1,
         N2919_1, N2921_1, N2922_1, N2934_1, N2935_1, N2936_1, N2937_1,
         N2979_1, N2981_1, N2982_1, N2994_1, N2995_1, N3023_1, N3024_1,
         N3025_1, N3026_1, N3401_1, N3402_1, N3403_1, N3404_1, N3409_1,
         N3410_1, N3411_1, N3412_1, N3445_1, N3446_1, N3450_1, N3451_1,
         N3452_1, N3459_1, N3460_1, N3461_1, N3462_1, N3481_1, N3483_1,
         N3484_1, N3489_1, N3490_1, N3504_1, N3505_1, N3506_1, N3507_1,
         N3616_1, N3617_1, N3618_1, N3619_1, N3620_1, N3621_1, N3622_1,
         N3623_1, N3624_1, N3627_1, N3628_1, N3629_1, N3630_1, N3631_1,
         N3632_1, N3633_1, N3634_1, N3635_1, N3638_1, N3641_1, N3642_1,
         N3643_1, N3644_1, N3645_1, N3646_1, N3647_1, N3648_1, N3649_1,
         N3650_1, N3651_1, N3652_1, N3653_1, N3654_1, N3655_1, N3656_1,
         N3657_1, N3658_1, N3659_1, N3660_1, N3661_1, N3662_1, N3663_1,
         N3668_1, N3669_1, N3670_1, N3671_1, N3676_1, N3677_1, N3678_1,
         N3679_1, N3703_1, N3704_1, N3711_1, N3712_1, N3713_1, N3719_1,
         N3720_1, N3721_1, N3722_1, N3745_1, N3746_1, N3747_1, N3751_1,
         N3752_1, N3758_1, N3760_1, N3767_1, N3768_1, N3769_1, N3770_1,
         N3781_1, N3782_1, N3783_1, N3784_1, N3785_1, N3786_1, N3787_1,
         N3788_1, N3800_1, N3801_1, N3802_1, N3803_1, N3804_1, N3805_1,
         N3806_1, N3807_1, N3808_1, N3809_1, N3980_1, N3981_1, N3998_1,
         N4032_1, N4033_1, N4034_1, N4035_1, N4037_1, N4038_1, N4039_1,
         N4040_1, N4185_1, N4186_1, N4196_1, N4197_1, N4273_1, N4273_2,
         N4274_1, N4274_2, N4276_1, N4276_2, N4277_1, N4277_2, N4547_1,
         N4741_1, N4953_1, N4954_1, N4955_1, N4956_1, N4957_1, N4958_1,
         N4959_1, N4960_1, N4961_1, N4978_1, N4979_1, N4980_1, N4981_1,
         N4982_1, N4983_1, N4984_1, N4985_1, N4986_1, N4987_1, N5060_1,
         N5060_2, N5061_1, N5061_2, N5062_1, N5062_2, N5063_1, N5063_2,
         N5066_1, N5068_1, N5163_1, N5164_1, N5165_1, N5240_1, N5388_1,
         N6072_1, N6073_1, N6073_2, N6074_1, N6074_2, N6076_1, N6077_1,
         N6077_2, N6078_1, N6078_2, N6080_1, N6080_2, N6084_1, N6085_1,
         N6087_1, N6091_1, N6091_2, N6091_3, N6095_1, N6096_1, N6096_2,
         N6097_1, N6097_2, N6097_3, N6099_1, N6100_1, N6100_2, N6101_1,
         N6101_2, N6101_3, N6103_1, N6104_1, N6104_2, N6106_1, N6108_1,
         N6108_2, N6112_1, N6113_1, N6115_1, N6117_1, N6117_2, N6117_3,
         N6121_1, N6122_1, N6122_2, N6123_1, N6123_2, N6123_3, N6125_1,
         N6126_1, N6126_2, N6127_1, N6127_2, N6129_1, N6130_1, N6130_2,
         N6132_1, N6133_1, N6135_1, N6140_1, N6140_2, N6143_1, N6144_1,
         N6145_1, N6149_1, N6149_2, N6149_3, N6153_1, N6154_1, N6154_2,
         N6155_1, N6155_2, N6155_3, N6156_1, N6157_1, N6157_2, N6158_1,
         N6158_2, N6158_3, N6160_1, N6161_1, N6161_2, N6163_1, N6168_1,
         N6168_2, N6171_1, N6172_1, N6173_1, N6175_1, N6175_2, N6175_3,
         N6179_1, N6180_1, N6180_2, N6181_1, N6181_2, N6181_3, N6182_1,
         N6183_1, N6183_2, N6184_1, N6184_2, N6185_1, N6186_1, N6186_2,
         N6188_1, N6189_1, N6191_1, N6382_1, N6382_2, N6386_1, N6386_2,
         N6388_1, N6388_2, N6392_1, N6392_2, N6397_1, N6397_2, N6397_3,
         N6415_1, N6415_2, N6415_3, N6427_1, N6427_2, N6427_3, N6441_1,
         N6441_2, N6441_3, N6473_1, N6474_1, N6475_1, N6476_1, N6482_1,
         N6482_2, N6490_1, N6500_1, N6500_2, N6500_3, N6504_1, N6504_2,
         N6508_1, N6516_1, N6516_2, N6536_1, N6536_2, N6539_1, N6539_2,
         N6539_3, N6556_1, N6556_2, N6566_1, N6566_2, N6572_1, N6580_1,
         N6580_2, N6580_3, N6584_1, N6584_2, N6587_1, N6592_1, N6592_2,
         N6606_1, N6606_2, N6609_1, N6609_2, N6609_3, N6622_1, N6622_2,
         N6712_1, N6713_1, N6714_1, N6715_1, N6718_1, N6719_1, N6720_1,
         N6721_1, N6722_1, N6860_1, N6861_1, N6862_1, N6863_1, N6866_1,
         N7011_1, N7012_1, N7013_1, N7016_1, N7114_1, N7146_1, N7147_1,
         N7187_1, N7188_1, N7189_1, N7190_1, N7196_1, N7197_1, N7198_1,
         N7207_1, N7208_1, N7270_1, N7276_1, N7282_1, N7288_1, N7294_1,
         N7304_1, N7310_1, N7338_1, N7339_1, N7340_1, N7341_1, N7342_1,
         N7349_1, N7357_1, N7364_1, N7433_1, N7434_1, N7435_1, N7435_2,
         N7436_1, N7437_1, N7438_1, N7439_1, N7440_1, N7441_1, N7442_1,
         N7443_1, N7443_2, N7444_1, N7445_1, N7446_1, N7447_1, N7448_1,
         N7449_1, N7449_2, N7450_1, N7451_1, N7452_1, N7453_1, N7454_1,
         N7455_1, N7456_1, N7457_1, N7458_1, N7459_1, N7460_1, N7461_1,
         N7462_1, N7463_1, N7464_1, N7469_1, N7469_2, N7481_1, N7482_1,
         N7483_1, N7484_1, N7485_1, N7486_1, N7487_1, N7488_1, N7503_1,
         N7503_2, N7503_3, N7503_4, N7503_5, N7503_6, N7503_7, N7504_1,
         N7504_2, N7504_3, N7504_4, N7504_5, N7504_6, N7504_7, N7505_1,
         N7505_2, N7507_1, N7507_2, N7508_1, N7508_2, N7509_1, N7509_2,
         N7510_1, N7510_2, N7512_1, N7512_2, N7513_1, N7513_2, N7514_1,
         N7514_2, N7515_1, N7515_2, N7516_1, N7516_2, N7517_1, N7517_2,
         N7518_1, N7518_2, N7519_1, N7519_2, N7520_1, N7520_2, N7521_1,
         N7521_2, N7522_1, N7522_2, N7525_1, N7525_2, N7526_1, N7531_1,
         N7537_1, N7543_1, N7549_1, N7555_1, N7561_1, N7567_1, N7573_1,
         N7631_1, N7631_2, N7631_3, N7636_1, N7666_1, N7667_1, N7668_1,
         N7669_1, N7670_1, N7671_1, N7672_1, N7673_1, N7674_1, N7675_1,
         N7676_1, N7677_1, N7678_1, N7679_1, N7680_1, N7681_1, N7682_1,
         N7683_1, N7684_1, N7685_1, N7686_1, N7687_1, N7688_1, N7689_1,
         N7690_1, N7691_1, N7692_1, N7693_1, N7694_1, N7695_1, N7696_1,
         N7697_1, N7703_1, N7727_1, N7727_2, N7728_1, N7728_2, N7729_1,
         N7729_2, N7730_1, N7730_2, N7731_1, N7731_2, N7732_1, N7732_2,
         N7733_1, N7733_2, N7734_1, N7734_2, N7735_1, N7735_2, N7736_1,
         N7736_2, N7737_1, N7737_2, N7738_1, N7738_2, N7739_1, N7739_2,
         N7740_1, N7740_2, N7741_1, N7741_2, N7742_1, N7742_2, N7988_1,
         N7989_1, N7990_1, N7991_1, N7994_1, N7995_1, N7996_1, N7997_1,
         N8013_1, N8013_2, N8017_1, N8017_2, N8071_1, N8072_1, N8075_1,
         N8075_2, N8076_1, N8076_2, N8113_1, N8114_1, N8115_1, N8116_1,
         N8117_1, N8118_1, N8119_1, N8120_1, N8121_1, N8121_2, N8122_1,
         N8122_2, N8123_1, N8123_2, N8124_1, N8124_2;

  BUFX2 gate1 ( .A(N141), .Y(N709) );
  BUFX2 gate2 ( .A(N293), .Y(N816) );
  AND2X1 gate3 ( .A(N135), .B(N631), .Y(N1042) );
  INVX1 gate4 ( .A(N591), .Y(N1043) );
  BUFX2 gate5 ( .A(N592), .Y(N1066) );
  INVX1 gate6 ( .A(N595), .Y(N1067) );
  INVX1 gate7 ( .A(N596), .Y(N1080) );
  INVX1 gate8 ( .A(N597), .Y(N1092) );
  INVX1 gate9 ( .A(N598), .Y(N1104) );
  INVX1 gate10 ( .A(N545), .Y(N1137) );
  INVX1 gate11 ( .A(N348), .Y(N1138) );
  INVX1 gate12 ( .A(N366), .Y(N1139) );
  AND2X1 gate13 ( .A(N552), .B(N562), .Y(N1140) );
  INVX1 gate14 ( .A(N549), .Y(N1141) );
  INVX1 gate15 ( .A(N545), .Y(N1142) );
  INVX1 gate16 ( .A(N545), .Y(N1143) );
  INVX1 gate17 ( .A(N338), .Y(N1144) );
  INVX1 gate18 ( .A(N358), .Y(N1145) );
  NAND2X1 gate19 ( .A(N373), .B(N1), .Y(N1146) );
  AND2X1 gate20 ( .A(N141), .B(N145), .Y(N1147) );
  INVX1 gate21 ( .A(N592), .Y(N1148) );
  INVX1 gate22 ( .A(N1042), .Y(N1149) );
  AND2X1 gate23 ( .A(N1043), .B(N27), .Y(N1150) );
  AND2X1 gate24 ( .A(N386), .B(N556), .Y(N1151) );
  INVX1 gate25 ( .A(N245), .Y(N1152) );
  INVX1 gate26 ( .A(N552), .Y(N1153) );
  INVX1 gate27 ( .A(N562), .Y(N1154) );
  INVX1 gate28 ( .A(N559), .Y(N1155) );
  AND2X1 gate29_1 ( .A(N386), .B(N559), .Y(N1156_1) );
  AND2X1 gate29_2 ( .A(N556), .B(N552), .Y(N1156_2) );
  AND2X1 gate29 ( .A(N1156_1), .B(N1156_2), .Y(N1156) );
  INVX1 gate30 ( .A(N566), .Y(N1157) );
  BUFX2 gate31 ( .A(N571), .Y(N1161) );
  BUFX2 gate32 ( .A(N574), .Y(N1173) );
  BUFX2 gate33 ( .A(N571), .Y(N1185) );
  BUFX2 gate34 ( .A(N574), .Y(N1197) );
  BUFX2 gate35 ( .A(N137), .Y(N1209) );
  BUFX2 gate36 ( .A(N137), .Y(N1213) );
  BUFX2 gate37 ( .A(N141), .Y(N1216) );
  INVX1 gate38 ( .A(N583), .Y(N1219) );
  BUFX2 gate39 ( .A(N577), .Y(N1223) );
  BUFX2 gate40 ( .A(N580), .Y(N1235) );
  BUFX2 gate41 ( .A(N577), .Y(N1247) );
  BUFX2 gate42 ( .A(N580), .Y(N1259) );
  BUFX2 gate43 ( .A(N254), .Y(N1271) );
  BUFX2 gate44 ( .A(N251), .Y(N1280) );
  BUFX2 gate45 ( .A(N251), .Y(N1292) );
  BUFX2 gate46 ( .A(N248), .Y(N1303) );
  BUFX2 gate47 ( .A(N248), .Y(N1315) );
  BUFX2 gate48 ( .A(N610), .Y(N1327) );
  BUFX2 gate49 ( .A(N607), .Y(N1339) );
  BUFX2 gate50 ( .A(N613), .Y(N1351) );
  BUFX2 gate51 ( .A(N616), .Y(N1363) );
  BUFX2 gate52 ( .A(N210), .Y(N1375) );
  BUFX2 gate53 ( .A(N210), .Y(N1378) );
  BUFX2 gate54 ( .A(N218), .Y(N1381) );
  BUFX2 gate55 ( .A(N218), .Y(N1384) );
  BUFX2 gate56 ( .A(N226), .Y(N1387) );
  BUFX2 gate57 ( .A(N226), .Y(N1390) );
  BUFX2 gate58 ( .A(N234), .Y(N1393) );
  BUFX2 gate59 ( .A(N234), .Y(N1396) );
  BUFX2 gate60 ( .A(N257), .Y(N1415) );
  BUFX2 gate61 ( .A(N257), .Y(N1418) );
  BUFX2 gate62 ( .A(N265), .Y(N1421) );
  BUFX2 gate63 ( .A(N265), .Y(N1424) );
  BUFX2 gate64 ( .A(N273), .Y(N1427) );
  BUFX2 gate65 ( .A(N273), .Y(N1430) );
  BUFX2 gate66 ( .A(N281), .Y(N1433) );
  BUFX2 gate67 ( .A(N281), .Y(N1436) );
  BUFX2 gate68 ( .A(N335), .Y(N1455) );
  BUFX2 gate69 ( .A(N335), .Y(N1462) );
  BUFX2 gate70 ( .A(N206), .Y(N1469) );
  AND2X1 gate71 ( .A(N27), .B(N31), .Y(N1475) );
  BUFX2 gate72 ( .A(N1), .Y(N1479) );
  BUFX2 gate73 ( .A(N588), .Y(N1482) );
  BUFX2 gate74 ( .A(N293), .Y(N1492) );
  BUFX2 gate75 ( .A(N302), .Y(N1495) );
  BUFX2 gate76 ( .A(N308), .Y(N1498) );
  BUFX2 gate77 ( .A(N308), .Y(N1501) );
  BUFX2 gate78 ( .A(N316), .Y(N1504) );
  BUFX2 gate79 ( .A(N316), .Y(N1507) );
  BUFX2 gate80 ( .A(N324), .Y(N1510) );
  BUFX2 gate81 ( .A(N324), .Y(N1513) );
  BUFX2 gate82 ( .A(N341), .Y(N1516) );
  BUFX2 gate83 ( .A(N341), .Y(N1519) );
  BUFX2 gate84 ( .A(N351), .Y(N1522) );
  BUFX2 gate85 ( .A(N351), .Y(N1525) );
  BUFX2 gate86 ( .A(N257), .Y(N1542) );
  BUFX2 gate87 ( .A(N257), .Y(N1545) );
  BUFX2 gate88 ( .A(N265), .Y(N1548) );
  BUFX2 gate89 ( .A(N265), .Y(N1551) );
  BUFX2 gate90 ( .A(N273), .Y(N1554) );
  BUFX2 gate91 ( .A(N273), .Y(N1557) );
  BUFX2 gate92 ( .A(N281), .Y(N1560) );
  BUFX2 gate93 ( .A(N281), .Y(N1563) );
  BUFX2 gate94 ( .A(N332), .Y(N1566) );
  BUFX2 gate95 ( .A(N332), .Y(N1573) );
  BUFX2 gate96 ( .A(N549), .Y(N1580) );
  AND2X1 gate97 ( .A(N31), .B(N27), .Y(N1583) );
  INVX1 gate98 ( .A(N588), .Y(N1588) );
  BUFX2 gate99 ( .A(N324), .Y(N1594) );
  BUFX2 gate100 ( .A(N324), .Y(N1597) );
  BUFX2 gate101 ( .A(N341), .Y(N1600) );
  BUFX2 gate102 ( .A(N341), .Y(N1603) );
  BUFX2 gate103 ( .A(N351), .Y(N1606) );
  BUFX2 gate104 ( .A(N351), .Y(N1609) );
  BUFX2 gate105 ( .A(N293), .Y(N1612) );
  BUFX2 gate106 ( .A(N302), .Y(N1615) );
  BUFX2 gate107 ( .A(N308), .Y(N1618) );
  BUFX2 gate108 ( .A(N308), .Y(N1621) );
  BUFX2 gate109 ( .A(N316), .Y(N1624) );
  BUFX2 gate110 ( .A(N316), .Y(N1627) );
  BUFX2 gate111 ( .A(N361), .Y(N1630) );
  BUFX2 gate112 ( .A(N361), .Y(N1633) );
  BUFX2 gate113 ( .A(N210), .Y(N1636) );
  BUFX2 gate114 ( .A(N210), .Y(N1639) );
  BUFX2 gate115 ( .A(N218), .Y(N1642) );
  BUFX2 gate116 ( .A(N218), .Y(N1645) );
  BUFX2 gate117 ( .A(N226), .Y(N1648) );
  BUFX2 gate118 ( .A(N226), .Y(N1651) );
  BUFX2 gate119 ( .A(N234), .Y(N1654) );
  BUFX2 gate120 ( .A(N234), .Y(N1657) );
  INVX1 gate121 ( .A(N324), .Y(N1660) );
  BUFX2 gate122 ( .A(N242), .Y(N1663) );
  BUFX2 gate123 ( .A(N242), .Y(N1675) );
  BUFX2 gate124 ( .A(N254), .Y(N1685) );
  BUFX2 gate125 ( .A(N610), .Y(N1697) );
  BUFX2 gate126 ( .A(N607), .Y(N1709) );
  BUFX2 gate127 ( .A(N625), .Y(N1721) );
  BUFX2 gate128 ( .A(N619), .Y(N1727) );
  BUFX2 gate129 ( .A(N613), .Y(N1731) );
  BUFX2 gate130 ( .A(N616), .Y(N1743) );
  INVX1 gate131 ( .A(N599), .Y(N1755) );
  INVX1 gate132 ( .A(N603), .Y(N1758) );
  BUFX2 gate133 ( .A(N619), .Y(N1761) );
  BUFX2 gate134 ( .A(N625), .Y(N1769) );
  BUFX2 gate135 ( .A(N619), .Y(N1777) );
  BUFX2 gate136 ( .A(N625), .Y(N1785) );
  BUFX2 gate137 ( .A(N619), .Y(N1793) );
  BUFX2 gate138 ( .A(N625), .Y(N1800) );
  BUFX2 gate139 ( .A(N619), .Y(N1807) );
  BUFX2 gate140 ( .A(N625), .Y(N1814) );
  BUFX2 gate141 ( .A(N299), .Y(N1821) );
  BUFX2 gate142 ( .A(N446), .Y(N1824) );
  BUFX2 gate143 ( .A(N457), .Y(N1827) );
  BUFX2 gate144 ( .A(N468), .Y(N1830) );
  BUFX2 gate145 ( .A(N422), .Y(N1833) );
  BUFX2 gate146 ( .A(N435), .Y(N1836) );
  BUFX2 gate147 ( .A(N389), .Y(N1839) );
  BUFX2 gate148 ( .A(N400), .Y(N1842) );
  BUFX2 gate149 ( .A(N411), .Y(N1845) );
  BUFX2 gate150 ( .A(N374), .Y(N1848) );
  BUFX2 gate151 ( .A(N4), .Y(N1851) );
  BUFX2 gate152 ( .A(N446), .Y(N1854) );
  BUFX2 gate153 ( .A(N457), .Y(N1857) );
  BUFX2 gate154 ( .A(N468), .Y(N1860) );
  BUFX2 gate155 ( .A(N435), .Y(N1863) );
  BUFX2 gate156 ( .A(N389), .Y(N1866) );
  BUFX2 gate157 ( .A(N400), .Y(N1869) );
  BUFX2 gate158 ( .A(N411), .Y(N1872) );
  BUFX2 gate159 ( .A(N422), .Y(N1875) );
  BUFX2 gate160 ( .A(N374), .Y(N1878) );
  BUFX2 gate161 ( .A(N479), .Y(N1881) );
  BUFX2 gate162 ( .A(N490), .Y(N1884) );
  BUFX2 gate163 ( .A(N503), .Y(N1887) );
  BUFX2 gate164 ( .A(N514), .Y(N1890) );
  BUFX2 gate165 ( .A(N523), .Y(N1893) );
  BUFX2 gate166 ( .A(N534), .Y(N1896) );
  BUFX2 gate167 ( .A(N54), .Y(N1899) );
  BUFX2 gate168 ( .A(N479), .Y(N1902) );
  BUFX2 gate169 ( .A(N503), .Y(N1905) );
  BUFX2 gate170 ( .A(N514), .Y(N1908) );
  BUFX2 gate171 ( .A(N523), .Y(N1911) );
  BUFX2 gate172 ( .A(N534), .Y(N1914) );
  BUFX2 gate173 ( .A(N490), .Y(N1917) );
  BUFX2 gate174 ( .A(N361), .Y(N1920) );
  BUFX2 gate175 ( .A(N369), .Y(N1923) );
  BUFX2 gate176 ( .A(N341), .Y(N1926) );
  BUFX2 gate177 ( .A(N351), .Y(N1929) );
  BUFX2 gate178 ( .A(N308), .Y(N1932) );
  BUFX2 gate179 ( .A(N316), .Y(N1935) );
  BUFX2 gate180 ( .A(N293), .Y(N1938) );
  BUFX2 gate181 ( .A(N302), .Y(N1941) );
  BUFX2 gate182 ( .A(N281), .Y(N1944) );
  BUFX2 gate183 ( .A(N289), .Y(N1947) );
  BUFX2 gate184 ( .A(N265), .Y(N1950) );
  BUFX2 gate185 ( .A(N273), .Y(N1953) );
  BUFX2 gate186 ( .A(N234), .Y(N1956) );
  BUFX2 gate187 ( .A(N257), .Y(N1959) );
  BUFX2 gate188 ( .A(N218), .Y(N1962) );
  BUFX2 gate189 ( .A(N226), .Y(N1965) );
  BUFX2 gate190 ( .A(N210), .Y(N1968) );
  INVX1 gate191 ( .A(N1146), .Y(N1972) );
  AND2X1 gate192 ( .A(N136), .B(N1148), .Y(N2054) );
  INVX1 gate193 ( .A(N1150), .Y(N2060) );
  INVX1 gate194 ( .A(N1151), .Y(N2061) );
  BUFX2 gate195 ( .A(N1209), .Y(N2139) );
  BUFX2 gate196 ( .A(N1216), .Y(N2142) );
  BUFX2 gate197 ( .A(N1479), .Y(N2309) );
  AND2X1 gate198 ( .A(N1104), .B(N514), .Y(N2349) );
  OR2X1 gate199 ( .A(N1067), .B(N514), .Y(N2350) );
  BUFX2 gate200 ( .A(N1580), .Y(N2387) );
  BUFX2 gate201 ( .A(N1821), .Y(N2527) );
  INVX1 gate202 ( .A(N1580), .Y(N2584) );
  AND2X1 gate203_1 ( .A(N170), .B(N1161), .Y(N2585_1) );
  AND2X1 gate203 ( .A(N1173), .B(N2585_1), .Y(N2585) );
  AND2X1 gate204_1 ( .A(N173), .B(N1161), .Y(N2586_1) );
  AND2X1 gate204 ( .A(N1173), .B(N2586_1), .Y(N2586) );
  AND2X1 gate205_1 ( .A(N167), .B(N1161), .Y(N2587_1) );
  AND2X1 gate205 ( .A(N1173), .B(N2587_1), .Y(N2587) );
  AND2X1 gate206_1 ( .A(N164), .B(N1161), .Y(N2588_1) );
  AND2X1 gate206 ( .A(N1173), .B(N2588_1), .Y(N2588) );
  AND2X1 gate207_1 ( .A(N161), .B(N1161), .Y(N2589_1) );
  AND2X1 gate207 ( .A(N1173), .B(N2589_1), .Y(N2589) );
  NAND2X1 gate208 ( .A(N1475), .B(N140), .Y(N2590) );
  AND2X1 gate209_1 ( .A(N185), .B(N1185), .Y(N2591_1) );
  AND2X1 gate209 ( .A(N1197), .B(N2591_1), .Y(N2591) );
  AND2X1 gate210_1 ( .A(N158), .B(N1185), .Y(N2592_1) );
  AND2X1 gate210 ( .A(N1197), .B(N2592_1), .Y(N2592) );
  AND2X1 gate211_1 ( .A(N152), .B(N1185), .Y(N2593_1) );
  AND2X1 gate211 ( .A(N1197), .B(N2593_1), .Y(N2593) );
  AND2X1 gate212_1 ( .A(N146), .B(N1185), .Y(N2594_1) );
  AND2X1 gate212 ( .A(N1197), .B(N2594_1), .Y(N2594) );
  AND2X1 gate213_1 ( .A(N170), .B(N1223), .Y(N2595_1) );
  AND2X1 gate213 ( .A(N1235), .B(N2595_1), .Y(N2595) );
  AND2X1 gate214_1 ( .A(N173), .B(N1223), .Y(N2596_1) );
  AND2X1 gate214 ( .A(N1235), .B(N2596_1), .Y(N2596) );
  AND2X1 gate215_1 ( .A(N167), .B(N1223), .Y(N2597_1) );
  AND2X1 gate215 ( .A(N1235), .B(N2597_1), .Y(N2597) );
  AND2X1 gate216_1 ( .A(N164), .B(N1223), .Y(N2598_1) );
  AND2X1 gate216 ( .A(N1235), .B(N2598_1), .Y(N2598) );
  AND2X1 gate217_1 ( .A(N161), .B(N1223), .Y(N2599_1) );
  AND2X1 gate217 ( .A(N1235), .B(N2599_1), .Y(N2599) );
  AND2X1 gate218_1 ( .A(N185), .B(N1247), .Y(N2600_1) );
  AND2X1 gate218 ( .A(N1259), .B(N2600_1), .Y(N2600) );
  AND2X1 gate219_1 ( .A(N158), .B(N1247), .Y(N2601_1) );
  AND2X1 gate219 ( .A(N1259), .B(N2601_1), .Y(N2601) );
  AND2X1 gate220_1 ( .A(N152), .B(N1247), .Y(N2602_1) );
  AND2X1 gate220 ( .A(N1259), .B(N2602_1), .Y(N2602) );
  AND2X1 gate221_1 ( .A(N146), .B(N1247), .Y(N2603_1) );
  AND2X1 gate221 ( .A(N1259), .B(N2603_1), .Y(N2603) );
  AND2X1 gate222_1 ( .A(N106), .B(N1731), .Y(N2604_1) );
  AND2X1 gate222 ( .A(N1743), .B(N2604_1), .Y(N2604) );
  AND2X1 gate223_1 ( .A(N61), .B(N1327), .Y(N2605_1) );
  AND2X1 gate223 ( .A(N1339), .B(N2605_1), .Y(N2605) );
  AND2X1 gate224_1 ( .A(N106), .B(N1697), .Y(N2606_1) );
  AND2X1 gate224 ( .A(N1709), .B(N2606_1), .Y(N2606) );
  AND2X1 gate225_1 ( .A(N49), .B(N1697), .Y(N2607_1) );
  AND2X1 gate225 ( .A(N1709), .B(N2607_1), .Y(N2607) );
  AND2X1 gate226_1 ( .A(N103), .B(N1697), .Y(N2608_1) );
  AND2X1 gate226 ( .A(N1709), .B(N2608_1), .Y(N2608) );
  AND2X1 gate227_1 ( .A(N40), .B(N1697), .Y(N2609_1) );
  AND2X1 gate227 ( .A(N1709), .B(N2609_1), .Y(N2609) );
  AND2X1 gate228_1 ( .A(N37), .B(N1697), .Y(N2610_1) );
  AND2X1 gate228 ( .A(N1709), .B(N2610_1), .Y(N2610) );
  AND2X1 gate229_1 ( .A(N20), .B(N1327), .Y(N2611_1) );
  AND2X1 gate229 ( .A(N1339), .B(N2611_1), .Y(N2611) );
  AND2X1 gate230_1 ( .A(N17), .B(N1327), .Y(N2612_1) );
  AND2X1 gate230 ( .A(N1339), .B(N2612_1), .Y(N2612) );
  AND2X1 gate231_1 ( .A(N70), .B(N1327), .Y(N2613_1) );
  AND2X1 gate231 ( .A(N1339), .B(N2613_1), .Y(N2613) );
  AND2X1 gate232_1 ( .A(N64), .B(N1327), .Y(N2614_1) );
  AND2X1 gate232 ( .A(N1339), .B(N2614_1), .Y(N2614) );
  AND2X1 gate233_1 ( .A(N49), .B(N1731), .Y(N2615_1) );
  AND2X1 gate233 ( .A(N1743), .B(N2615_1), .Y(N2615) );
  AND2X1 gate234_1 ( .A(N103), .B(N1731), .Y(N2616_1) );
  AND2X1 gate234 ( .A(N1743), .B(N2616_1), .Y(N2616) );
  AND2X1 gate235_1 ( .A(N40), .B(N1731), .Y(N2617_1) );
  AND2X1 gate235 ( .A(N1743), .B(N2617_1), .Y(N2617) );
  AND2X1 gate236_1 ( .A(N37), .B(N1731), .Y(N2618_1) );
  AND2X1 gate236 ( .A(N1743), .B(N2618_1), .Y(N2618) );
  AND2X1 gate237_1 ( .A(N20), .B(N1351), .Y(N2619_1) );
  AND2X1 gate237 ( .A(N1363), .B(N2619_1), .Y(N2619) );
  AND2X1 gate238_1 ( .A(N17), .B(N1351), .Y(N2620_1) );
  AND2X1 gate238 ( .A(N1363), .B(N2620_1), .Y(N2620) );
  AND2X1 gate239_1 ( .A(N70), .B(N1351), .Y(N2621_1) );
  AND2X1 gate239 ( .A(N1363), .B(N2621_1), .Y(N2621) );
  AND2X1 gate240_1 ( .A(N64), .B(N1351), .Y(N2622_1) );
  AND2X1 gate240 ( .A(N1363), .B(N2622_1), .Y(N2622) );
  INVX1 gate241 ( .A(N1475), .Y(N2623) );
  AND2X1 gate242_1 ( .A(N123), .B(N1758), .Y(N2624_1) );
  AND2X1 gate242 ( .A(N599), .B(N2624_1), .Y(N2624) );
  AND2X1 gate243 ( .A(N1777), .B(N1785), .Y(N2625) );
  AND2X1 gate244_1 ( .A(N61), .B(N1351), .Y(N2626_1) );
  AND2X1 gate244 ( .A(N1363), .B(N2626_1), .Y(N2626) );
  AND2X1 gate245 ( .A(N1761), .B(N1769), .Y(N2627) );
  INVX1 gate246 ( .A(N1824), .Y(N2628) );
  INVX1 gate247 ( .A(N1827), .Y(N2629) );
  INVX1 gate248 ( .A(N1830), .Y(N2630) );
  INVX1 gate249 ( .A(N1833), .Y(N2631) );
  INVX1 gate250 ( .A(N1836), .Y(N2632) );
  INVX1 gate251 ( .A(N1839), .Y(N2633) );
  INVX1 gate252 ( .A(N1842), .Y(N2634) );
  INVX1 gate253 ( .A(N1845), .Y(N2635) );
  INVX1 gate254 ( .A(N1848), .Y(N2636) );
  INVX1 gate255 ( .A(N1851), .Y(N2637) );
  INVX1 gate256 ( .A(N1854), .Y(N2638) );
  INVX1 gate257 ( .A(N1857), .Y(N2639) );
  INVX1 gate258 ( .A(N1860), .Y(N2640) );
  INVX1 gate259 ( .A(N1863), .Y(N2641) );
  INVX1 gate260 ( .A(N1866), .Y(N2642) );
  INVX1 gate261 ( .A(N1869), .Y(N2643) );
  INVX1 gate262 ( .A(N1872), .Y(N2644) );
  INVX1 gate263 ( .A(N1875), .Y(N2645) );
  INVX1 gate264 ( .A(N1878), .Y(N2646) );
  BUFX2 gate265 ( .A(N1209), .Y(N2647) );
  INVX1 gate266 ( .A(N1161), .Y(N2653) );
  INVX1 gate267 ( .A(N1173), .Y(N2664) );
  BUFX2 gate268 ( .A(N1209), .Y(N2675) );
  INVX1 gate269 ( .A(N1185), .Y(N2681) );
  INVX1 gate270 ( .A(N1197), .Y(N2692) );
  AND2X1 gate271_1 ( .A(N179), .B(N1185), .Y(N2703_1) );
  AND2X1 gate271 ( .A(N1197), .B(N2703_1), .Y(N2703) );
  BUFX2 gate272 ( .A(N1479), .Y(N2704) );
  INVX1 gate273 ( .A(N1881), .Y(N2709) );
  INVX1 gate274 ( .A(N1884), .Y(N2710) );
  INVX1 gate275 ( .A(N1887), .Y(N2711) );
  INVX1 gate276 ( .A(N1890), .Y(N2712) );
  INVX1 gate277 ( .A(N1893), .Y(N2713) );
  INVX1 gate278 ( .A(N1896), .Y(N2714) );
  INVX1 gate279 ( .A(N1899), .Y(N2715) );
  INVX1 gate280 ( .A(N1902), .Y(N2716) );
  INVX1 gate281 ( .A(N1905), .Y(N2717) );
  INVX1 gate282 ( .A(N1908), .Y(N2718) );
  INVX1 gate283 ( .A(N1911), .Y(N2719) );
  INVX1 gate284 ( .A(N1914), .Y(N2720) );
  INVX1 gate285 ( .A(N1917), .Y(N2721) );
  BUFX2 gate286 ( .A(N1213), .Y(N2722) );
  INVX1 gate287 ( .A(N1223), .Y(N2728) );
  INVX1 gate288 ( .A(N1235), .Y(N2739) );
  BUFX2 gate289 ( .A(N1213), .Y(N2750) );
  INVX1 gate290 ( .A(N1247), .Y(N2756) );
  INVX1 gate291 ( .A(N1259), .Y(N2767) );
  AND2X1 gate292_1 ( .A(N179), .B(N1247), .Y(N2778_1) );
  AND2X1 gate292 ( .A(N1259), .B(N2778_1), .Y(N2778) );
  INVX1 gate293 ( .A(N1327), .Y(N2779) );
  INVX1 gate294 ( .A(N1339), .Y(N2790) );
  INVX1 gate295 ( .A(N1351), .Y(N2801) );
  INVX1 gate296 ( .A(N1363), .Y(N2812) );
  INVX1 gate297 ( .A(N1375), .Y(N2823) );
  INVX1 gate298 ( .A(N1378), .Y(N2824) );
  INVX1 gate299 ( .A(N1381), .Y(N2825) );
  INVX1 gate300 ( .A(N1384), .Y(N2826) );
  INVX1 gate301 ( .A(N1387), .Y(N2827) );
  INVX1 gate302 ( .A(N1390), .Y(N2828) );
  INVX1 gate303 ( .A(N1393), .Y(N2829) );
  INVX1 gate304 ( .A(N1396), .Y(N2830) );
  AND2X1 gate305_1 ( .A(N1104), .B(N457), .Y(N2831_1) );
  AND2X1 gate305 ( .A(N1378), .B(N2831_1), .Y(N2831) );
  AND2X1 gate306_1 ( .A(N1104), .B(N468), .Y(N2832_1) );
  AND2X1 gate306 ( .A(N1384), .B(N2832_1), .Y(N2832) );
  AND2X1 gate307_1 ( .A(N1104), .B(N422), .Y(N2833_1) );
  AND2X1 gate307 ( .A(N1390), .B(N2833_1), .Y(N2833) );
  AND2X1 gate308_1 ( .A(N1104), .B(N435), .Y(N2834_1) );
  AND2X1 gate308 ( .A(N1396), .B(N2834_1), .Y(N2834) );
  AND2X1 gate309 ( .A(N1067), .B(N1375), .Y(N2835) );
  AND2X1 gate310 ( .A(N1067), .B(N1381), .Y(N2836) );
  AND2X1 gate311 ( .A(N1067), .B(N1387), .Y(N2837) );
  AND2X1 gate312 ( .A(N1067), .B(N1393), .Y(N2838) );
  INVX1 gate313 ( .A(N1415), .Y(N2839) );
  INVX1 gate314 ( .A(N1418), .Y(N2840) );
  INVX1 gate315 ( .A(N1421), .Y(N2841) );
  INVX1 gate316 ( .A(N1424), .Y(N2842) );
  INVX1 gate317 ( .A(N1427), .Y(N2843) );
  INVX1 gate318 ( .A(N1430), .Y(N2844) );
  INVX1 gate319 ( .A(N1433), .Y(N2845) );
  INVX1 gate320 ( .A(N1436), .Y(N2846) );
  AND2X1 gate321_1 ( .A(N1104), .B(N389), .Y(N2847_1) );
  AND2X1 gate321 ( .A(N1418), .B(N2847_1), .Y(N2847) );
  AND2X1 gate322_1 ( .A(N1104), .B(N400), .Y(N2848_1) );
  AND2X1 gate322 ( .A(N1424), .B(N2848_1), .Y(N2848) );
  AND2X1 gate323_1 ( .A(N1104), .B(N411), .Y(N2849_1) );
  AND2X1 gate323 ( .A(N1430), .B(N2849_1), .Y(N2849) );
  AND2X1 gate324_1 ( .A(N1104), .B(N374), .Y(N2850_1) );
  AND2X1 gate324 ( .A(N1436), .B(N2850_1), .Y(N2850) );
  AND2X1 gate325 ( .A(N1067), .B(N1415), .Y(N2851) );
  AND2X1 gate326 ( .A(N1067), .B(N1421), .Y(N2852) );
  AND2X1 gate327 ( .A(N1067), .B(N1427), .Y(N2853) );
  AND2X1 gate328 ( .A(N1067), .B(N1433), .Y(N2854) );
  INVX1 gate329 ( .A(N1455), .Y(N2855) );
  INVX1 gate330 ( .A(N1462), .Y(N2861) );
  AND2X1 gate331 ( .A(N292), .B(N1455), .Y(N2867) );
  AND2X1 gate332 ( .A(N288), .B(N1455), .Y(N2868) );
  AND2X1 gate333 ( .A(N280), .B(N1455), .Y(N2869) );
  AND2X1 gate334 ( .A(N272), .B(N1455), .Y(N2870) );
  AND2X1 gate335 ( .A(N264), .B(N1455), .Y(N2871) );
  AND2X1 gate336 ( .A(N241), .B(N1462), .Y(N2872) );
  AND2X1 gate337 ( .A(N233), .B(N1462), .Y(N2873) );
  AND2X1 gate338 ( .A(N225), .B(N1462), .Y(N2874) );
  AND2X1 gate339 ( .A(N217), .B(N1462), .Y(N2875) );
  AND2X1 gate340 ( .A(N209), .B(N1462), .Y(N2876) );
  BUFX2 gate341 ( .A(N1216), .Y(N2877) );
  INVX1 gate342 ( .A(N1482), .Y(N2882) );
  INVX1 gate343 ( .A(N1475), .Y(N2891) );
  INVX1 gate344 ( .A(N1492), .Y(N2901) );
  INVX1 gate345 ( .A(N1495), .Y(N2902) );
  INVX1 gate346 ( .A(N1498), .Y(N2903) );
  INVX1 gate347 ( .A(N1501), .Y(N2904) );
  INVX1 gate348 ( .A(N1504), .Y(N2905) );
  INVX1 gate349 ( .A(N1507), .Y(N2906) );
  AND2X1 gate350 ( .A(N1303), .B(N1495), .Y(N2907) );
  AND2X1 gate351_1 ( .A(N1303), .B(N479), .Y(N2908_1) );
  AND2X1 gate351 ( .A(N1501), .B(N2908_1), .Y(N2908) );
  AND2X1 gate352_1 ( .A(N1303), .B(N490), .Y(N2909_1) );
  AND2X1 gate352 ( .A(N1507), .B(N2909_1), .Y(N2909) );
  AND2X1 gate353 ( .A(N1663), .B(N1492), .Y(N2910) );
  AND2X1 gate354 ( .A(N1663), .B(N1498), .Y(N2911) );
  AND2X1 gate355 ( .A(N1663), .B(N1504), .Y(N2912) );
  INVX1 gate356 ( .A(N1510), .Y(N2913) );
  INVX1 gate357 ( .A(N1513), .Y(N2914) );
  INVX1 gate358 ( .A(N1516), .Y(N2915) );
  INVX1 gate359 ( .A(N1519), .Y(N2916) );
  INVX1 gate360 ( .A(N1522), .Y(N2917) );
  INVX1 gate361 ( .A(N1525), .Y(N2918) );
  AND2X1 gate362_1 ( .A(N1104), .B(N503), .Y(N2919_1) );
  AND2X1 gate362 ( .A(N1513), .B(N2919_1), .Y(N2919) );
  INVX1 gate363 ( .A(N2349), .Y(N2920) );
  AND2X1 gate364_1 ( .A(N1104), .B(N523), .Y(N2921_1) );
  AND2X1 gate364 ( .A(N1519), .B(N2921_1), .Y(N2921) );
  AND2X1 gate365_1 ( .A(N1104), .B(N534), .Y(N2922_1) );
  AND2X1 gate365 ( .A(N1525), .B(N2922_1), .Y(N2922) );
  AND2X1 gate366 ( .A(N1067), .B(N1510), .Y(N2923) );
  AND2X1 gate367 ( .A(N1067), .B(N1516), .Y(N2924) );
  AND2X1 gate368 ( .A(N1067), .B(N1522), .Y(N2925) );
  INVX1 gate369 ( .A(N1542), .Y(N2926) );
  INVX1 gate370 ( .A(N1545), .Y(N2927) );
  INVX1 gate371 ( .A(N1548), .Y(N2928) );
  INVX1 gate372 ( .A(N1551), .Y(N2929) );
  INVX1 gate373 ( .A(N1554), .Y(N2930) );
  INVX1 gate374 ( .A(N1557), .Y(N2931) );
  INVX1 gate375 ( .A(N1560), .Y(N2932) );
  INVX1 gate376 ( .A(N1563), .Y(N2933) );
  AND2X1 gate377_1 ( .A(N1303), .B(N389), .Y(N2934_1) );
  AND2X1 gate377 ( .A(N1545), .B(N2934_1), .Y(N2934) );
  AND2X1 gate378_1 ( .A(N1303), .B(N400), .Y(N2935_1) );
  AND2X1 gate378 ( .A(N1551), .B(N2935_1), .Y(N2935) );
  AND2X1 gate379_1 ( .A(N1303), .B(N411), .Y(N2936_1) );
  AND2X1 gate379 ( .A(N1557), .B(N2936_1), .Y(N2936) );
  AND2X1 gate380_1 ( .A(N1303), .B(N374), .Y(N2937_1) );
  AND2X1 gate380 ( .A(N1563), .B(N2937_1), .Y(N2937) );
  AND2X1 gate381 ( .A(N1663), .B(N1542), .Y(N2938) );
  AND2X1 gate382 ( .A(N1663), .B(N1548), .Y(N2939) );
  AND2X1 gate383 ( .A(N1663), .B(N1554), .Y(N2940) );
  AND2X1 gate384 ( .A(N1663), .B(N1560), .Y(N2941) );
  INVX1 gate385 ( .A(N1566), .Y(N2942) );
  INVX1 gate386 ( .A(N1573), .Y(N2948) );
  AND2X1 gate387 ( .A(N372), .B(N1566), .Y(N2954) );
  AND2X1 gate388 ( .A(N366), .B(N1566), .Y(N2955) );
  AND2X1 gate389 ( .A(N358), .B(N1566), .Y(N2956) );
  AND2X1 gate390 ( .A(N348), .B(N1566), .Y(N2957) );
  AND2X1 gate391 ( .A(N338), .B(N1566), .Y(N2958) );
  AND2X1 gate392 ( .A(N331), .B(N1573), .Y(N2959) );
  AND2X1 gate393 ( .A(N323), .B(N1573), .Y(N2960) );
  AND2X1 gate394 ( .A(N315), .B(N1573), .Y(N2961) );
  AND2X1 gate395 ( .A(N307), .B(N1573), .Y(N2962) );
  AND2X1 gate396 ( .A(N299), .B(N1573), .Y(N2963) );
  INVX1 gate397 ( .A(N1588), .Y(N2964) );
  AND2X1 gate398 ( .A(N83), .B(N1588), .Y(N2969) );
  AND2X1 gate399 ( .A(N86), .B(N1588), .Y(N2970) );
  AND2X1 gate400 ( .A(N88), .B(N1588), .Y(N2971) );
  AND2X1 gate401 ( .A(N88), .B(N1588), .Y(N2972) );
  INVX1 gate402 ( .A(N1594), .Y(N2973) );
  INVX1 gate403 ( .A(N1597), .Y(N2974) );
  INVX1 gate404 ( .A(N1600), .Y(N2975) );
  INVX1 gate405 ( .A(N1603), .Y(N2976) );
  INVX1 gate406 ( .A(N1606), .Y(N2977) );
  INVX1 gate407 ( .A(N1609), .Y(N2978) );
  AND2X1 gate408_1 ( .A(N1315), .B(N503), .Y(N2979_1) );
  AND2X1 gate408 ( .A(N1597), .B(N2979_1), .Y(N2979) );
  AND2X1 gate409 ( .A(N1315), .B(N514), .Y(N2980) );
  AND2X1 gate410_1 ( .A(N1315), .B(N523), .Y(N2981_1) );
  AND2X1 gate410 ( .A(N1603), .B(N2981_1), .Y(N2981) );
  AND2X1 gate411_1 ( .A(N1315), .B(N534), .Y(N2982_1) );
  AND2X1 gate411 ( .A(N1609), .B(N2982_1), .Y(N2982) );
  AND2X1 gate412 ( .A(N1675), .B(N1594), .Y(N2983) );
  OR2X1 gate413 ( .A(N1675), .B(N514), .Y(N2984) );
  AND2X1 gate414 ( .A(N1675), .B(N1600), .Y(N2985) );
  AND2X1 gate415 ( .A(N1675), .B(N1606), .Y(N2986) );
  INVX1 gate416 ( .A(N1612), .Y(N2987) );
  INVX1 gate417 ( .A(N1615), .Y(N2988) );
  INVX1 gate418 ( .A(N1618), .Y(N2989) );
  INVX1 gate419 ( .A(N1621), .Y(N2990) );
  INVX1 gate420 ( .A(N1624), .Y(N2991) );
  INVX1 gate421 ( .A(N1627), .Y(N2992) );
  AND2X1 gate422 ( .A(N1315), .B(N1615), .Y(N2993) );
  AND2X1 gate423_1 ( .A(N1315), .B(N479), .Y(N2994_1) );
  AND2X1 gate423 ( .A(N1621), .B(N2994_1), .Y(N2994) );
  AND2X1 gate424_1 ( .A(N1315), .B(N490), .Y(N2995_1) );
  AND2X1 gate424 ( .A(N1627), .B(N2995_1), .Y(N2995) );
  AND2X1 gate425 ( .A(N1675), .B(N1612), .Y(N2996) );
  AND2X1 gate426 ( .A(N1675), .B(N1618), .Y(N2997) );
  AND2X1 gate427 ( .A(N1675), .B(N1624), .Y(N2998) );
  INVX1 gate428 ( .A(N1630), .Y(N2999) );
  BUFX2 gate429 ( .A(N1469), .Y(N3000) );
  BUFX2 gate430 ( .A(N1469), .Y(N3003) );
  INVX1 gate431 ( .A(N1633), .Y(N3006) );
  BUFX2 gate432 ( .A(N1469), .Y(N3007) );
  BUFX2 gate433 ( .A(N1469), .Y(N3010) );
  AND2X1 gate434 ( .A(N1315), .B(N1630), .Y(N3013) );
  AND2X1 gate435 ( .A(N1315), .B(N1633), .Y(N3014) );
  INVX1 gate436 ( .A(N1636), .Y(N3015) );
  INVX1 gate437 ( .A(N1639), .Y(N3016) );
  INVX1 gate438 ( .A(N1642), .Y(N3017) );
  INVX1 gate439 ( .A(N1645), .Y(N3018) );
  INVX1 gate440 ( .A(N1648), .Y(N3019) );
  INVX1 gate441 ( .A(N1651), .Y(N3020) );
  INVX1 gate442 ( .A(N1654), .Y(N3021) );
  INVX1 gate443 ( .A(N1657), .Y(N3022) );
  AND2X1 gate444_1 ( .A(N1303), .B(N457), .Y(N3023_1) );
  AND2X1 gate444 ( .A(N1639), .B(N3023_1), .Y(N3023) );
  AND2X1 gate445_1 ( .A(N1303), .B(N468), .Y(N3024_1) );
  AND2X1 gate445 ( .A(N1645), .B(N3024_1), .Y(N3024) );
  AND2X1 gate446_1 ( .A(N1303), .B(N422), .Y(N3025_1) );
  AND2X1 gate446 ( .A(N1651), .B(N3025_1), .Y(N3025) );
  AND2X1 gate447_1 ( .A(N1303), .B(N435), .Y(N3026_1) );
  AND2X1 gate447 ( .A(N1657), .B(N3026_1), .Y(N3026) );
  AND2X1 gate448 ( .A(N1663), .B(N1636), .Y(N3027) );
  AND2X1 gate449 ( .A(N1663), .B(N1642), .Y(N3028) );
  AND2X1 gate450 ( .A(N1663), .B(N1648), .Y(N3029) );
  AND2X1 gate451 ( .A(N1663), .B(N1654), .Y(N3030) );
  INVX1 gate452 ( .A(N1920), .Y(N3031) );
  INVX1 gate453 ( .A(N1923), .Y(N3032) );
  INVX1 gate454 ( .A(N1926), .Y(N3033) );
  INVX1 gate455 ( .A(N1929), .Y(N3034) );
  BUFX2 gate456 ( .A(N1660), .Y(N3035) );
  BUFX2 gate457 ( .A(N1660), .Y(N3038) );
  INVX1 gate458 ( .A(N1697), .Y(N3041) );
  INVX1 gate459 ( .A(N1709), .Y(N3052) );
  INVX1 gate460 ( .A(N1721), .Y(N3063) );
  INVX1 gate461 ( .A(N1727), .Y(N3068) );
  AND2X1 gate462 ( .A(N97), .B(N1721), .Y(N3071) );
  AND2X1 gate463 ( .A(N94), .B(N1721), .Y(N3072) );
  AND2X1 gate464 ( .A(N97), .B(N1721), .Y(N3073) );
  AND2X1 gate465 ( .A(N94), .B(N1721), .Y(N3074) );
  INVX1 gate466 ( .A(N1731), .Y(N3075) );
  INVX1 gate467 ( .A(N1743), .Y(N3086) );
  INVX1 gate468 ( .A(N1761), .Y(N3097) );
  INVX1 gate469 ( .A(N1769), .Y(N3108) );
  INVX1 gate470 ( .A(N1777), .Y(N3119) );
  INVX1 gate471 ( .A(N1785), .Y(N3130) );
  INVX1 gate472 ( .A(N1944), .Y(N3141) );
  INVX1 gate473 ( .A(N1947), .Y(N3142) );
  INVX1 gate474 ( .A(N1950), .Y(N3143) );
  INVX1 gate475 ( .A(N1953), .Y(N3144) );
  INVX1 gate476 ( .A(N1956), .Y(N3145) );
  INVX1 gate477 ( .A(N1959), .Y(N3146) );
  INVX1 gate478 ( .A(N1793), .Y(N3147) );
  INVX1 gate479 ( .A(N1800), .Y(N3158) );
  INVX1 gate480 ( .A(N1807), .Y(N3169) );
  INVX1 gate481 ( .A(N1814), .Y(N3180) );
  BUFX2 gate482 ( .A(N1821), .Y(N3191) );
  INVX1 gate483 ( .A(N1932), .Y(N3194) );
  INVX1 gate484 ( .A(N1935), .Y(N3195) );
  INVX1 gate485 ( .A(N1938), .Y(N3196) );
  INVX1 gate486 ( .A(N1941), .Y(N3197) );
  INVX1 gate487 ( .A(N1962), .Y(N3198) );
  INVX1 gate488 ( .A(N1965), .Y(N3199) );
  BUFX2 gate489 ( .A(N1469), .Y(N3200) );
  INVX1 gate490 ( .A(N1968), .Y(N3203) );
  BUFX2 gate491 ( .A(N2704), .Y(N3357) );
  BUFX2 gate492 ( .A(N2704), .Y(N3358) );
  BUFX2 gate493 ( .A(N2704), .Y(N3359) );
  BUFX2 gate494 ( .A(N2704), .Y(N3360) );
  AND2X1 gate495_1 ( .A(N457), .B(N1092), .Y(N3401_1) );
  AND2X1 gate495 ( .A(N2824), .B(N3401_1), .Y(N3401) );
  AND2X1 gate496_1 ( .A(N468), .B(N1092), .Y(N3402_1) );
  AND2X1 gate496 ( .A(N2826), .B(N3402_1), .Y(N3402) );
  AND2X1 gate497_1 ( .A(N422), .B(N1092), .Y(N3403_1) );
  AND2X1 gate497 ( .A(N2828), .B(N3403_1), .Y(N3403) );
  AND2X1 gate498_1 ( .A(N435), .B(N1092), .Y(N3404_1) );
  AND2X1 gate498 ( .A(N2830), .B(N3404_1), .Y(N3404) );
  AND2X1 gate499 ( .A(N1080), .B(N2823), .Y(N3405) );
  AND2X1 gate500 ( .A(N1080), .B(N2825), .Y(N3406) );
  AND2X1 gate501 ( .A(N1080), .B(N2827), .Y(N3407) );
  AND2X1 gate502 ( .A(N1080), .B(N2829), .Y(N3408) );
  AND2X1 gate503_1 ( .A(N389), .B(N1092), .Y(N3409_1) );
  AND2X1 gate503 ( .A(N2840), .B(N3409_1), .Y(N3409) );
  AND2X1 gate504_1 ( .A(N400), .B(N1092), .Y(N3410_1) );
  AND2X1 gate504 ( .A(N2842), .B(N3410_1), .Y(N3410) );
  AND2X1 gate505_1 ( .A(N411), .B(N1092), .Y(N3411_1) );
  AND2X1 gate505 ( .A(N2844), .B(N3411_1), .Y(N3411) );
  AND2X1 gate506_1 ( .A(N374), .B(N1092), .Y(N3412_1) );
  AND2X1 gate506 ( .A(N2846), .B(N3412_1), .Y(N3412) );
  AND2X1 gate507 ( .A(N1080), .B(N2839), .Y(N3413) );
  AND2X1 gate508 ( .A(N1080), .B(N2841), .Y(N3414) );
  AND2X1 gate509 ( .A(N1080), .B(N2843), .Y(N3415) );
  AND2X1 gate510 ( .A(N1080), .B(N2845), .Y(N3416) );
  AND2X1 gate511 ( .A(N1280), .B(N2902), .Y(N3444) );
  AND2X1 gate512_1 ( .A(N479), .B(N1280), .Y(N3445_1) );
  AND2X1 gate512 ( .A(N2904), .B(N3445_1), .Y(N3445) );
  AND2X1 gate513_1 ( .A(N490), .B(N1280), .Y(N3446_1) );
  AND2X1 gate513 ( .A(N2906), .B(N3446_1), .Y(N3446) );
  AND2X1 gate514 ( .A(N1685), .B(N2901), .Y(N3447) );
  AND2X1 gate515 ( .A(N1685), .B(N2903), .Y(N3448) );
  AND2X1 gate516 ( .A(N1685), .B(N2905), .Y(N3449) );
  AND2X1 gate517_1 ( .A(N503), .B(N1092), .Y(N3450_1) );
  AND2X1 gate517 ( .A(N2914), .B(N3450_1), .Y(N3450) );
  AND2X1 gate518_1 ( .A(N523), .B(N1092), .Y(N3451_1) );
  AND2X1 gate518 ( .A(N2916), .B(N3451_1), .Y(N3451) );
  AND2X1 gate519_1 ( .A(N534), .B(N1092), .Y(N3452_1) );
  AND2X1 gate519 ( .A(N2918), .B(N3452_1), .Y(N3452) );
  AND2X1 gate520 ( .A(N1080), .B(N2913), .Y(N3453) );
  AND2X1 gate521 ( .A(N1080), .B(N2915), .Y(N3454) );
  AND2X1 gate522 ( .A(N1080), .B(N2917), .Y(N3455) );
  AND2X1 gate523 ( .A(N2920), .B(N2350), .Y(N3456) );
  AND2X1 gate524_1 ( .A(N389), .B(N1280), .Y(N3459_1) );
  AND2X1 gate524 ( .A(N2927), .B(N3459_1), .Y(N3459) );
  AND2X1 gate525_1 ( .A(N400), .B(N1280), .Y(N3460_1) );
  AND2X1 gate525 ( .A(N2929), .B(N3460_1), .Y(N3460) );
  AND2X1 gate526_1 ( .A(N411), .B(N1280), .Y(N3461_1) );
  AND2X1 gate526 ( .A(N2931), .B(N3461_1), .Y(N3461) );
  AND2X1 gate527_1 ( .A(N374), .B(N1280), .Y(N3462_1) );
  AND2X1 gate527 ( .A(N2933), .B(N3462_1), .Y(N3462) );
  AND2X1 gate528 ( .A(N1685), .B(N2926), .Y(N3463) );
  AND2X1 gate529 ( .A(N1685), .B(N2928), .Y(N3464) );
  AND2X1 gate530 ( .A(N1685), .B(N2930), .Y(N3465) );
  AND2X1 gate531 ( .A(N1685), .B(N2932), .Y(N3466) );
  AND2X1 gate532_1 ( .A(N503), .B(N1292), .Y(N3481_1) );
  AND2X1 gate532 ( .A(N2974), .B(N3481_1), .Y(N3481) );
  INVX1 gate533 ( .A(N2980), .Y(N3482) );
  AND2X1 gate534_1 ( .A(N523), .B(N1292), .Y(N3483_1) );
  AND2X1 gate534 ( .A(N2976), .B(N3483_1), .Y(N3483) );
  AND2X1 gate535_1 ( .A(N534), .B(N1292), .Y(N3484_1) );
  AND2X1 gate535 ( .A(N2978), .B(N3484_1), .Y(N3484) );
  AND2X1 gate536 ( .A(N1271), .B(N2973), .Y(N3485) );
  AND2X1 gate537 ( .A(N1271), .B(N2975), .Y(N3486) );
  AND2X1 gate538 ( .A(N1271), .B(N2977), .Y(N3487) );
  AND2X1 gate539 ( .A(N1292), .B(N2988), .Y(N3488) );
  AND2X1 gate540_1 ( .A(N479), .B(N1292), .Y(N3489_1) );
  AND2X1 gate540 ( .A(N2990), .B(N3489_1), .Y(N3489) );
  AND2X1 gate541_1 ( .A(N490), .B(N1292), .Y(N3490_1) );
  AND2X1 gate541 ( .A(N2992), .B(N3490_1), .Y(N3490) );
  AND2X1 gate542 ( .A(N1271), .B(N2987), .Y(N3491) );
  AND2X1 gate543 ( .A(N1271), .B(N2989), .Y(N3492) );
  AND2X1 gate544 ( .A(N1271), .B(N2991), .Y(N3493) );
  AND2X1 gate545 ( .A(N1292), .B(N2999), .Y(N3502) );
  AND2X1 gate546 ( .A(N1292), .B(N3006), .Y(N3503) );
  AND2X1 gate547_1 ( .A(N457), .B(N1280), .Y(N3504_1) );
  AND2X1 gate547 ( .A(N3016), .B(N3504_1), .Y(N3504) );
  AND2X1 gate548_1 ( .A(N468), .B(N1280), .Y(N3505_1) );
  AND2X1 gate548 ( .A(N3018), .B(N3505_1), .Y(N3505) );
  AND2X1 gate549_1 ( .A(N422), .B(N1280), .Y(N3506_1) );
  AND2X1 gate549 ( .A(N3020), .B(N3506_1), .Y(N3506) );
  AND2X1 gate550_1 ( .A(N435), .B(N1280), .Y(N3507_1) );
  AND2X1 gate550 ( .A(N3022), .B(N3507_1), .Y(N3507) );
  AND2X1 gate551 ( .A(N1685), .B(N3015), .Y(N3508) );
  AND2X1 gate552 ( .A(N1685), .B(N3017), .Y(N3509) );
  AND2X1 gate553 ( .A(N1685), .B(N3019), .Y(N3510) );
  AND2X1 gate554 ( .A(N1685), .B(N3021), .Y(N3511) );
  NAND2X1 gate555 ( .A(N1923), .B(N3031), .Y(N3512) );
  NAND2X1 gate556 ( .A(N1920), .B(N3032), .Y(N3513) );
  NAND2X1 gate557 ( .A(N1929), .B(N3033), .Y(N3514) );
  NAND2X1 gate558 ( .A(N1926), .B(N3034), .Y(N3515) );
  NAND2X1 gate559 ( .A(N1947), .B(N3141), .Y(N3558) );
  NAND2X1 gate560 ( .A(N1944), .B(N3142), .Y(N3559) );
  NAND2X1 gate561 ( .A(N1953), .B(N3143), .Y(N3560) );
  NAND2X1 gate562 ( .A(N1950), .B(N3144), .Y(N3561) );
  NAND2X1 gate563 ( .A(N1959), .B(N3145), .Y(N3562) );
  NAND2X1 gate564 ( .A(N1956), .B(N3146), .Y(N3563) );
  BUFX2 gate565 ( .A(N3191), .Y(N3604) );
  NAND2X1 gate566 ( .A(N1935), .B(N3194), .Y(N3605) );
  NAND2X1 gate567 ( .A(N1932), .B(N3195), .Y(N3606) );
  NAND2X1 gate568 ( .A(N1941), .B(N3196), .Y(N3607) );
  NAND2X1 gate569 ( .A(N1938), .B(N3197), .Y(N3608) );
  NAND2X1 gate570 ( .A(N1965), .B(N3198), .Y(N3609) );
  NAND2X1 gate571 ( .A(N1962), .B(N3199), .Y(N3610) );
  INVX1 gate572 ( .A(N3191), .Y(N3613) );
  AND2X1 gate573 ( .A(N2882), .B(N2891), .Y(N3614) );
  AND2X1 gate574 ( .A(N1482), .B(N2891), .Y(N3615) );
  AND2X1 gate575_1 ( .A(N200), .B(N2653), .Y(N3616_1) );
  AND2X1 gate575 ( .A(N1173), .B(N3616_1), .Y(N3616) );
  AND2X1 gate576_1 ( .A(N203), .B(N2653), .Y(N3617_1) );
  AND2X1 gate576 ( .A(N1173), .B(N3617_1), .Y(N3617) );
  AND2X1 gate577_1 ( .A(N197), .B(N2653), .Y(N3618_1) );
  AND2X1 gate577 ( .A(N1173), .B(N3618_1), .Y(N3618) );
  AND2X1 gate578_1 ( .A(N194), .B(N2653), .Y(N3619_1) );
  AND2X1 gate578 ( .A(N1173), .B(N3619_1), .Y(N3619) );
  AND2X1 gate579_1 ( .A(N191), .B(N2653), .Y(N3620_1) );
  AND2X1 gate579 ( .A(N1173), .B(N3620_1), .Y(N3620) );
  AND2X1 gate580_1 ( .A(N182), .B(N2681), .Y(N3621_1) );
  AND2X1 gate580 ( .A(N1197), .B(N3621_1), .Y(N3621) );
  AND2X1 gate581_1 ( .A(N188), .B(N2681), .Y(N3622_1) );
  AND2X1 gate581 ( .A(N1197), .B(N3622_1), .Y(N3622) );
  AND2X1 gate582_1 ( .A(N155), .B(N2681), .Y(N3623_1) );
  AND2X1 gate582 ( .A(N1197), .B(N3623_1), .Y(N3623) );
  AND2X1 gate583_1 ( .A(N149), .B(N2681), .Y(N3624_1) );
  AND2X1 gate583 ( .A(N1197), .B(N3624_1), .Y(N3624) );
  AND2X1 gate584 ( .A(N2882), .B(N2891), .Y(N3625) );
  AND2X1 gate585 ( .A(N1482), .B(N2891), .Y(N3626) );
  AND2X1 gate586_1 ( .A(N200), .B(N2728), .Y(N3627_1) );
  AND2X1 gate586 ( .A(N1235), .B(N3627_1), .Y(N3627) );
  AND2X1 gate587_1 ( .A(N203), .B(N2728), .Y(N3628_1) );
  AND2X1 gate587 ( .A(N1235), .B(N3628_1), .Y(N3628) );
  AND2X1 gate588_1 ( .A(N197), .B(N2728), .Y(N3629_1) );
  AND2X1 gate588 ( .A(N1235), .B(N3629_1), .Y(N3629) );
  AND2X1 gate589_1 ( .A(N194), .B(N2728), .Y(N3630_1) );
  AND2X1 gate589 ( .A(N1235), .B(N3630_1), .Y(N3630) );
  AND2X1 gate590_1 ( .A(N191), .B(N2728), .Y(N3631_1) );
  AND2X1 gate590 ( .A(N1235), .B(N3631_1), .Y(N3631) );
  AND2X1 gate591_1 ( .A(N182), .B(N2756), .Y(N3632_1) );
  AND2X1 gate591 ( .A(N1259), .B(N3632_1), .Y(N3632) );
  AND2X1 gate592_1 ( .A(N188), .B(N2756), .Y(N3633_1) );
  AND2X1 gate592 ( .A(N1259), .B(N3633_1), .Y(N3633) );
  AND2X1 gate593_1 ( .A(N155), .B(N2756), .Y(N3634_1) );
  AND2X1 gate593 ( .A(N1259), .B(N3634_1), .Y(N3634) );
  AND2X1 gate594_1 ( .A(N149), .B(N2756), .Y(N3635_1) );
  AND2X1 gate594 ( .A(N1259), .B(N3635_1), .Y(N3635) );
  AND2X1 gate595 ( .A(N2882), .B(N2891), .Y(N3636) );
  AND2X1 gate596 ( .A(N1482), .B(N2891), .Y(N3637) );
  AND2X1 gate597_1 ( .A(N109), .B(N3075), .Y(N3638_1) );
  AND2X1 gate597 ( .A(N1743), .B(N3638_1), .Y(N3638) );
  AND2X1 gate598 ( .A(N2882), .B(N2891), .Y(N3639) );
  AND2X1 gate599 ( .A(N1482), .B(N2891), .Y(N3640) );
  AND2X1 gate600_1 ( .A(N11), .B(N2779), .Y(N3641_1) );
  AND2X1 gate600 ( .A(N1339), .B(N3641_1), .Y(N3641) );
  AND2X1 gate601_1 ( .A(N109), .B(N3041), .Y(N3642_1) );
  AND2X1 gate601 ( .A(N1709), .B(N3642_1), .Y(N3642) );
  AND2X1 gate602_1 ( .A(N46), .B(N3041), .Y(N3643_1) );
  AND2X1 gate602 ( .A(N1709), .B(N3643_1), .Y(N3643) );
  AND2X1 gate603_1 ( .A(N100), .B(N3041), .Y(N3644_1) );
  AND2X1 gate603 ( .A(N1709), .B(N3644_1), .Y(N3644) );
  AND2X1 gate604_1 ( .A(N91), .B(N3041), .Y(N3645_1) );
  AND2X1 gate604 ( .A(N1709), .B(N3645_1), .Y(N3645) );
  AND2X1 gate605_1 ( .A(N43), .B(N3041), .Y(N3646_1) );
  AND2X1 gate605 ( .A(N1709), .B(N3646_1), .Y(N3646) );
  AND2X1 gate606_1 ( .A(N76), .B(N2779), .Y(N3647_1) );
  AND2X1 gate606 ( .A(N1339), .B(N3647_1), .Y(N3647) );
  AND2X1 gate607_1 ( .A(N73), .B(N2779), .Y(N3648_1) );
  AND2X1 gate607 ( .A(N1339), .B(N3648_1), .Y(N3648) );
  AND2X1 gate608_1 ( .A(N67), .B(N2779), .Y(N3649_1) );
  AND2X1 gate608 ( .A(N1339), .B(N3649_1), .Y(N3649) );
  AND2X1 gate609_1 ( .A(N14), .B(N2779), .Y(N3650_1) );
  AND2X1 gate609 ( .A(N1339), .B(N3650_1), .Y(N3650) );
  AND2X1 gate610_1 ( .A(N46), .B(N3075), .Y(N3651_1) );
  AND2X1 gate610 ( .A(N1743), .B(N3651_1), .Y(N3651) );
  AND2X1 gate611_1 ( .A(N100), .B(N3075), .Y(N3652_1) );
  AND2X1 gate611 ( .A(N1743), .B(N3652_1), .Y(N3652) );
  AND2X1 gate612_1 ( .A(N91), .B(N3075), .Y(N3653_1) );
  AND2X1 gate612 ( .A(N1743), .B(N3653_1), .Y(N3653) );
  AND2X1 gate613_1 ( .A(N43), .B(N3075), .Y(N3654_1) );
  AND2X1 gate613 ( .A(N1743), .B(N3654_1), .Y(N3654) );
  AND2X1 gate614_1 ( .A(N76), .B(N2801), .Y(N3655_1) );
  AND2X1 gate614 ( .A(N1363), .B(N3655_1), .Y(N3655) );
  AND2X1 gate615_1 ( .A(N73), .B(N2801), .Y(N3656_1) );
  AND2X1 gate615 ( .A(N1363), .B(N3656_1), .Y(N3656) );
  AND2X1 gate616_1 ( .A(N67), .B(N2801), .Y(N3657_1) );
  AND2X1 gate616 ( .A(N1363), .B(N3657_1), .Y(N3657) );
  AND2X1 gate617_1 ( .A(N14), .B(N2801), .Y(N3658_1) );
  AND2X1 gate617 ( .A(N1363), .B(N3658_1), .Y(N3658) );
  AND2X1 gate618_1 ( .A(N120), .B(N3119), .Y(N3659_1) );
  AND2X1 gate618 ( .A(N1785), .B(N3659_1), .Y(N3659) );
  AND2X1 gate619_1 ( .A(N11), .B(N2801), .Y(N3660_1) );
  AND2X1 gate619 ( .A(N1363), .B(N3660_1), .Y(N3660) );
  AND2X1 gate620_1 ( .A(N118), .B(N3097), .Y(N3661_1) );
  AND2X1 gate620 ( .A(N1769), .B(N3661_1), .Y(N3661) );
  AND2X1 gate621_1 ( .A(N176), .B(N2681), .Y(N3662_1) );
  AND2X1 gate621 ( .A(N1197), .B(N3662_1), .Y(N3662) );
  AND2X1 gate622_1 ( .A(N176), .B(N2756), .Y(N3663_1) );
  AND2X1 gate622 ( .A(N1259), .B(N3663_1), .Y(N3663) );
  OR2X1 gate623 ( .A(N2831), .B(N3401), .Y(N3664) );
  OR2X1 gate624 ( .A(N2832), .B(N3402), .Y(N3665) );
  OR2X1 gate625 ( .A(N2833), .B(N3403), .Y(N3666) );
  OR2X1 gate626 ( .A(N2834), .B(N3404), .Y(N3667) );
  OR2X1 gate627_1 ( .A(N2835), .B(N3405), .Y(N3668_1) );
  OR2X1 gate627 ( .A(N457), .B(N3668_1), .Y(N3668) );
  OR2X1 gate628_1 ( .A(N2836), .B(N3406), .Y(N3669_1) );
  OR2X1 gate628 ( .A(N468), .B(N3669_1), .Y(N3669) );
  OR2X1 gate629_1 ( .A(N2837), .B(N3407), .Y(N3670_1) );
  OR2X1 gate629 ( .A(N422), .B(N3670_1), .Y(N3670) );
  OR2X1 gate630_1 ( .A(N2838), .B(N3408), .Y(N3671_1) );
  OR2X1 gate630 ( .A(N435), .B(N3671_1), .Y(N3671) );
  OR2X1 gate631 ( .A(N2847), .B(N3409), .Y(N3672) );
  OR2X1 gate632 ( .A(N2848), .B(N3410), .Y(N3673) );
  OR2X1 gate633 ( .A(N2849), .B(N3411), .Y(N3674) );
  OR2X1 gate634 ( .A(N2850), .B(N3412), .Y(N3675) );
  OR2X1 gate635_1 ( .A(N2851), .B(N3413), .Y(N3676_1) );
  OR2X1 gate635 ( .A(N389), .B(N3676_1), .Y(N3676) );
  OR2X1 gate636_1 ( .A(N2852), .B(N3414), .Y(N3677_1) );
  OR2X1 gate636 ( .A(N400), .B(N3677_1), .Y(N3677) );
  OR2X1 gate637_1 ( .A(N2853), .B(N3415), .Y(N3678_1) );
  OR2X1 gate637 ( .A(N411), .B(N3678_1), .Y(N3678) );
  OR2X1 gate638_1 ( .A(N2854), .B(N3416), .Y(N3679_1) );
  OR2X1 gate638 ( .A(N374), .B(N3679_1), .Y(N3679) );
  AND2X1 gate639 ( .A(N289), .B(N2855), .Y(N3680) );
  AND2X1 gate640 ( .A(N281), .B(N2855), .Y(N3681) );
  AND2X1 gate641 ( .A(N273), .B(N2855), .Y(N3682) );
  AND2X1 gate642 ( .A(N265), .B(N2855), .Y(N3683) );
  AND2X1 gate643 ( .A(N257), .B(N2855), .Y(N3684) );
  AND2X1 gate644 ( .A(N234), .B(N2861), .Y(N3685) );
  AND2X1 gate645 ( .A(N226), .B(N2861), .Y(N3686) );
  AND2X1 gate646 ( .A(N218), .B(N2861), .Y(N3687) );
  AND2X1 gate647 ( .A(N210), .B(N2861), .Y(N3688) );
  AND2X1 gate648 ( .A(N206), .B(N2861), .Y(N3689) );
  INVX1 gate649 ( .A(N2891), .Y(N3691) );
  OR2X1 gate650 ( .A(N2907), .B(N3444), .Y(N3700) );
  OR2X1 gate651 ( .A(N2908), .B(N3445), .Y(N3701) );
  OR2X1 gate652 ( .A(N2909), .B(N3446), .Y(N3702) );
  OR2X1 gate653_1 ( .A(N2911), .B(N3448), .Y(N3703_1) );
  OR2X1 gate653 ( .A(N479), .B(N3703_1), .Y(N3703) );
  OR2X1 gate654_1 ( .A(N2912), .B(N3449), .Y(N3704_1) );
  OR2X1 gate654 ( .A(N490), .B(N3704_1), .Y(N3704) );
  OR2X1 gate655 ( .A(N2910), .B(N3447), .Y(N3705) );
  OR2X1 gate656 ( .A(N2919), .B(N3450), .Y(N3708) );
  OR2X1 gate657 ( .A(N2921), .B(N3451), .Y(N3709) );
  OR2X1 gate658 ( .A(N2922), .B(N3452), .Y(N3710) );
  OR2X1 gate659_1 ( .A(N2923), .B(N3453), .Y(N3711_1) );
  OR2X1 gate659 ( .A(N503), .B(N3711_1), .Y(N3711) );
  OR2X1 gate660_1 ( .A(N2924), .B(N3454), .Y(N3712_1) );
  OR2X1 gate660 ( .A(N523), .B(N3712_1), .Y(N3712) );
  OR2X1 gate661_1 ( .A(N2925), .B(N3455), .Y(N3713_1) );
  OR2X1 gate661 ( .A(N534), .B(N3713_1), .Y(N3713) );
  OR2X1 gate662 ( .A(N2934), .B(N3459), .Y(N3715) );
  OR2X1 gate663 ( .A(N2935), .B(N3460), .Y(N3716) );
  OR2X1 gate664 ( .A(N2936), .B(N3461), .Y(N3717) );
  OR2X1 gate665 ( .A(N2937), .B(N3462), .Y(N3718) );
  OR2X1 gate666_1 ( .A(N2938), .B(N3463), .Y(N3719_1) );
  OR2X1 gate666 ( .A(N389), .B(N3719_1), .Y(N3719) );
  OR2X1 gate667_1 ( .A(N2939), .B(N3464), .Y(N3720_1) );
  OR2X1 gate667 ( .A(N400), .B(N3720_1), .Y(N3720) );
  OR2X1 gate668_1 ( .A(N2940), .B(N3465), .Y(N3721_1) );
  OR2X1 gate668 ( .A(N411), .B(N3721_1), .Y(N3721) );
  OR2X1 gate669_1 ( .A(N2941), .B(N3466), .Y(N3722_1) );
  OR2X1 gate669 ( .A(N374), .B(N3722_1), .Y(N3722) );
  AND2X1 gate670 ( .A(N369), .B(N2942), .Y(N3723) );
  AND2X1 gate671 ( .A(N361), .B(N2942), .Y(N3724) );
  AND2X1 gate672 ( .A(N351), .B(N2942), .Y(N3725) );
  AND2X1 gate673 ( .A(N341), .B(N2942), .Y(N3726) );
  AND2X1 gate674 ( .A(N324), .B(N2948), .Y(N3727) );
  AND2X1 gate675 ( .A(N316), .B(N2948), .Y(N3728) );
  AND2X1 gate676 ( .A(N308), .B(N2948), .Y(N3729) );
  AND2X1 gate677 ( .A(N302), .B(N2948), .Y(N3730) );
  AND2X1 gate678 ( .A(N293), .B(N2948), .Y(N3731) );
  OR2X1 gate679 ( .A(N2942), .B(N2958), .Y(N3732) );
  AND2X1 gate680 ( .A(N83), .B(N2964), .Y(N3738) );
  AND2X1 gate681 ( .A(N87), .B(N2964), .Y(N3739) );
  AND2X1 gate682 ( .A(N34), .B(N2964), .Y(N3740) );
  AND2X1 gate683 ( .A(N34), .B(N2964), .Y(N3741) );
  OR2X1 gate684 ( .A(N2979), .B(N3481), .Y(N3742) );
  OR2X1 gate685 ( .A(N2981), .B(N3483), .Y(N3743) );
  OR2X1 gate686 ( .A(N2982), .B(N3484), .Y(N3744) );
  OR2X1 gate687_1 ( .A(N2983), .B(N3485), .Y(N3745_1) );
  OR2X1 gate687 ( .A(N503), .B(N3745_1), .Y(N3745) );
  OR2X1 gate688_1 ( .A(N2985), .B(N3486), .Y(N3746_1) );
  OR2X1 gate688 ( .A(N523), .B(N3746_1), .Y(N3746) );
  OR2X1 gate689_1 ( .A(N2986), .B(N3487), .Y(N3747_1) );
  OR2X1 gate689 ( .A(N534), .B(N3747_1), .Y(N3747) );
  OR2X1 gate690 ( .A(N2993), .B(N3488), .Y(N3748) );
  OR2X1 gate691 ( .A(N2994), .B(N3489), .Y(N3749) );
  OR2X1 gate692 ( .A(N2995), .B(N3490), .Y(N3750) );
  OR2X1 gate693_1 ( .A(N2997), .B(N3492), .Y(N3751_1) );
  OR2X1 gate693 ( .A(N479), .B(N3751_1), .Y(N3751) );
  OR2X1 gate694_1 ( .A(N2998), .B(N3493), .Y(N3752_1) );
  OR2X1 gate694 ( .A(N490), .B(N3752_1), .Y(N3752) );
  INVX1 gate695 ( .A(N3000), .Y(N3753) );
  INVX1 gate696 ( .A(N3003), .Y(N3754) );
  INVX1 gate697 ( .A(N3007), .Y(N3755) );
  INVX1 gate698 ( .A(N3010), .Y(N3756) );
  OR2X1 gate699 ( .A(N3013), .B(N3502), .Y(N3757) );
  AND2X1 gate700_1 ( .A(N1315), .B(N446), .Y(N3758_1) );
  AND2X1 gate700 ( .A(N3003), .B(N3758_1), .Y(N3758) );
  OR2X1 gate701 ( .A(N3014), .B(N3503), .Y(N3759) );
  AND2X1 gate702_1 ( .A(N1315), .B(N446), .Y(N3760_1) );
  AND2X1 gate702 ( .A(N3010), .B(N3760_1), .Y(N3760) );
  AND2X1 gate703 ( .A(N1675), .B(N3000), .Y(N3761) );
  AND2X1 gate704 ( .A(N1675), .B(N3007), .Y(N3762) );
  OR2X1 gate705 ( .A(N3023), .B(N3504), .Y(N3763) );
  OR2X1 gate706 ( .A(N3024), .B(N3505), .Y(N3764) );
  OR2X1 gate707 ( .A(N3025), .B(N3506), .Y(N3765) );
  OR2X1 gate708 ( .A(N3026), .B(N3507), .Y(N3766) );
  OR2X1 gate709_1 ( .A(N3027), .B(N3508), .Y(N3767_1) );
  OR2X1 gate709 ( .A(N457), .B(N3767_1), .Y(N3767) );
  OR2X1 gate710_1 ( .A(N3028), .B(N3509), .Y(N3768_1) );
  OR2X1 gate710 ( .A(N468), .B(N3768_1), .Y(N3768) );
  OR2X1 gate711_1 ( .A(N3029), .B(N3510), .Y(N3769_1) );
  OR2X1 gate711 ( .A(N422), .B(N3769_1), .Y(N3769) );
  OR2X1 gate712_1 ( .A(N3030), .B(N3511), .Y(N3770_1) );
  OR2X1 gate712 ( .A(N435), .B(N3770_1), .Y(N3770) );
  NAND2X1 gate713 ( .A(N3512), .B(N3513), .Y(N3771) );
  NAND2X1 gate714 ( .A(N3514), .B(N3515), .Y(N3775) );
  INVX1 gate715 ( .A(N3035), .Y(N3779) );
  INVX1 gate716 ( .A(N3038), .Y(N3780) );
  AND2X1 gate717_1 ( .A(N117), .B(N3097), .Y(N3781_1) );
  AND2X1 gate717 ( .A(N1769), .B(N3781_1), .Y(N3781) );
  AND2X1 gate718_1 ( .A(N126), .B(N3097), .Y(N3782_1) );
  AND2X1 gate718 ( .A(N1769), .B(N3782_1), .Y(N3782) );
  AND2X1 gate719_1 ( .A(N127), .B(N3097), .Y(N3783_1) );
  AND2X1 gate719 ( .A(N1769), .B(N3783_1), .Y(N3783) );
  AND2X1 gate720_1 ( .A(N128), .B(N3097), .Y(N3784_1) );
  AND2X1 gate720 ( .A(N1769), .B(N3784_1), .Y(N3784) );
  AND2X1 gate721_1 ( .A(N131), .B(N3119), .Y(N3785_1) );
  AND2X1 gate721 ( .A(N1785), .B(N3785_1), .Y(N3785) );
  AND2X1 gate722_1 ( .A(N129), .B(N3119), .Y(N3786_1) );
  AND2X1 gate722 ( .A(N1785), .B(N3786_1), .Y(N3786) );
  AND2X1 gate723_1 ( .A(N119), .B(N3119), .Y(N3787_1) );
  AND2X1 gate723 ( .A(N1785), .B(N3787_1), .Y(N3787) );
  AND2X1 gate724_1 ( .A(N130), .B(N3119), .Y(N3788_1) );
  AND2X1 gate724 ( .A(N1785), .B(N3788_1), .Y(N3788) );
  NAND2X1 gate725 ( .A(N3558), .B(N3559), .Y(N3789) );
  NAND2X1 gate726 ( .A(N3560), .B(N3561), .Y(N3793) );
  NAND2X1 gate727 ( .A(N3562), .B(N3563), .Y(N3797) );
  AND2X1 gate728_1 ( .A(N122), .B(N3147), .Y(N3800_1) );
  AND2X1 gate728 ( .A(N1800), .B(N3800_1), .Y(N3800) );
  AND2X1 gate729_1 ( .A(N113), .B(N3147), .Y(N3801_1) );
  AND2X1 gate729 ( .A(N1800), .B(N3801_1), .Y(N3801) );
  AND2X1 gate730_1 ( .A(N53), .B(N3147), .Y(N3802_1) );
  AND2X1 gate730 ( .A(N1800), .B(N3802_1), .Y(N3802) );
  AND2X1 gate731_1 ( .A(N114), .B(N3147), .Y(N3803_1) );
  AND2X1 gate731 ( .A(N1800), .B(N3803_1), .Y(N3803) );
  AND2X1 gate732_1 ( .A(N115), .B(N3147), .Y(N3804_1) );
  AND2X1 gate732 ( .A(N1800), .B(N3804_1), .Y(N3804) );
  AND2X1 gate733_1 ( .A(N52), .B(N3169), .Y(N3805_1) );
  AND2X1 gate733 ( .A(N1814), .B(N3805_1), .Y(N3805) );
  AND2X1 gate734_1 ( .A(N112), .B(N3169), .Y(N3806_1) );
  AND2X1 gate734 ( .A(N1814), .B(N3806_1), .Y(N3806) );
  AND2X1 gate735_1 ( .A(N116), .B(N3169), .Y(N3807_1) );
  AND2X1 gate735 ( .A(N1814), .B(N3807_1), .Y(N3807) );
  AND2X1 gate736_1 ( .A(N121), .B(N3169), .Y(N3808_1) );
  AND2X1 gate736 ( .A(N1814), .B(N3808_1), .Y(N3808) );
  AND2X1 gate737_1 ( .A(N123), .B(N3169), .Y(N3809_1) );
  AND2X1 gate737 ( .A(N1814), .B(N3809_1), .Y(N3809) );
  NAND2X1 gate738 ( .A(N3607), .B(N3608), .Y(N3810) );
  NAND2X1 gate739 ( .A(N3605), .B(N3606), .Y(N3813) );
  AND2X1 gate740 ( .A(N3482), .B(N2984), .Y(N3816) );
  OR2X1 gate741 ( .A(N2996), .B(N3491), .Y(N3819) );
  INVX1 gate742 ( .A(N3200), .Y(N3822) );
  NAND2X1 gate743 ( .A(N3200), .B(N3203), .Y(N3823) );
  NAND2X1 gate744 ( .A(N3609), .B(N3610), .Y(N3824) );
  INVX1 gate745 ( .A(N3456), .Y(N3827) );
  OR2X1 gate746 ( .A(N3739), .B(N2970), .Y(N3828) );
  OR2X1 gate747 ( .A(N3740), .B(N2971), .Y(N3829) );
  OR2X1 gate748 ( .A(N3741), .B(N2972), .Y(N3830) );
  OR2X1 gate749 ( .A(N3738), .B(N2969), .Y(N3831) );
  INVX1 gate750 ( .A(N3664), .Y(N3834) );
  INVX1 gate751 ( .A(N3665), .Y(N3835) );
  INVX1 gate752 ( .A(N3666), .Y(N3836) );
  INVX1 gate753 ( .A(N3667), .Y(N3837) );
  INVX1 gate754 ( .A(N3672), .Y(N3838) );
  INVX1 gate755 ( .A(N3673), .Y(N3839) );
  INVX1 gate756 ( .A(N3674), .Y(N3840) );
  INVX1 gate757 ( .A(N3675), .Y(N3841) );
  OR2X1 gate758 ( .A(N3681), .B(N2868), .Y(N3842) );
  OR2X1 gate759 ( .A(N3682), .B(N2869), .Y(N3849) );
  OR2X1 gate760 ( .A(N3683), .B(N2870), .Y(N3855) );
  OR2X1 gate761 ( .A(N3684), .B(N2871), .Y(N3861) );
  OR2X1 gate762 ( .A(N3685), .B(N2872), .Y(N3867) );
  OR2X1 gate763 ( .A(N3686), .B(N2873), .Y(N3873) );
  OR2X1 gate764 ( .A(N3687), .B(N2874), .Y(N3881) );
  OR2X1 gate765 ( .A(N3688), .B(N2875), .Y(N3887) );
  OR2X1 gate766 ( .A(N3689), .B(N2876), .Y(N3893) );
  INVX1 gate767 ( .A(N3701), .Y(N3908) );
  INVX1 gate768 ( .A(N3702), .Y(N3909) );
  INVX1 gate769 ( .A(N3700), .Y(N3911) );
  INVX1 gate770 ( .A(N3708), .Y(N3914) );
  INVX1 gate771 ( .A(N3709), .Y(N3915) );
  INVX1 gate772 ( .A(N3710), .Y(N3916) );
  INVX1 gate773 ( .A(N3715), .Y(N3917) );
  INVX1 gate774 ( .A(N3716), .Y(N3918) );
  INVX1 gate775 ( .A(N3717), .Y(N3919) );
  INVX1 gate776 ( .A(N3718), .Y(N3920) );
  OR2X1 gate777 ( .A(N3724), .B(N2955), .Y(N3921) );
  OR2X1 gate778 ( .A(N3725), .B(N2956), .Y(N3927) );
  OR2X1 gate779 ( .A(N3726), .B(N2957), .Y(N3933) );
  OR2X1 gate780 ( .A(N3727), .B(N2959), .Y(N3942) );
  OR2X1 gate781 ( .A(N3728), .B(N2960), .Y(N3948) );
  OR2X1 gate782 ( .A(N3729), .B(N2961), .Y(N3956) );
  OR2X1 gate783 ( .A(N3730), .B(N2962), .Y(N3962) );
  OR2X1 gate784 ( .A(N3731), .B(N2963), .Y(N3968) );
  INVX1 gate785 ( .A(N3742), .Y(N3975) );
  INVX1 gate786 ( .A(N3743), .Y(N3976) );
  INVX1 gate787 ( .A(N3744), .Y(N3977) );
  INVX1 gate788 ( .A(N3749), .Y(N3978) );
  INVX1 gate789 ( .A(N3750), .Y(N3979) );
  AND2X1 gate790_1 ( .A(N446), .B(N1292), .Y(N3980_1) );
  AND2X1 gate790 ( .A(N3754), .B(N3980_1), .Y(N3980) );
  AND2X1 gate791_1 ( .A(N446), .B(N1292), .Y(N3981_1) );
  AND2X1 gate791 ( .A(N3756), .B(N3981_1), .Y(N3981) );
  AND2X1 gate792 ( .A(N1271), .B(N3753), .Y(N3982) );
  AND2X1 gate793 ( .A(N1271), .B(N3755), .Y(N3983) );
  INVX1 gate794 ( .A(N3757), .Y(N3984) );
  INVX1 gate795 ( .A(N3759), .Y(N3987) );
  INVX1 gate796 ( .A(N3763), .Y(N3988) );
  INVX1 gate797 ( .A(N3764), .Y(N3989) );
  INVX1 gate798 ( .A(N3765), .Y(N3990) );
  INVX1 gate799 ( .A(N3766), .Y(N3991) );
  AND2X1 gate800_1 ( .A(N3456), .B(N3119), .Y(N3998_1) );
  AND2X1 gate800 ( .A(N3130), .B(N3998_1), .Y(N3998) );
  OR2X1 gate801 ( .A(N3723), .B(N2954), .Y(N4008) );
  OR2X1 gate802 ( .A(N3680), .B(N2867), .Y(N4011) );
  INVX1 gate803 ( .A(N3748), .Y(N4021) );
  NAND2X1 gate804 ( .A(N1968), .B(N3822), .Y(N4024) );
  INVX1 gate805 ( .A(N3705), .Y(N4027) );
  AND2X1 gate806 ( .A(N3828), .B(N1583), .Y(N4031) );
  AND2X1 gate807_1 ( .A(N24), .B(N2882), .Y(N4032_1) );
  AND2X1 gate807 ( .A(N3691), .B(N4032_1), .Y(N4032) );
  AND2X1 gate808_1 ( .A(N25), .B(N1482), .Y(N4033_1) );
  AND2X1 gate808 ( .A(N3691), .B(N4033_1), .Y(N4033) );
  AND2X1 gate809_1 ( .A(N26), .B(N2882), .Y(N4034_1) );
  AND2X1 gate809 ( .A(N3691), .B(N4034_1), .Y(N4034) );
  AND2X1 gate810_1 ( .A(N81), .B(N1482), .Y(N4035_1) );
  AND2X1 gate810 ( .A(N3691), .B(N4035_1), .Y(N4035) );
  AND2X1 gate811 ( .A(N3829), .B(N1583), .Y(N4036) );
  AND2X1 gate812_1 ( .A(N79), .B(N2882), .Y(N4037_1) );
  AND2X1 gate812 ( .A(N3691), .B(N4037_1), .Y(N4037) );
  AND2X1 gate813_1 ( .A(N23), .B(N1482), .Y(N4038_1) );
  AND2X1 gate813 ( .A(N3691), .B(N4038_1), .Y(N4038) );
  AND2X1 gate814_1 ( .A(N82), .B(N2882), .Y(N4039_1) );
  AND2X1 gate814 ( .A(N3691), .B(N4039_1), .Y(N4039) );
  AND2X1 gate815_1 ( .A(N80), .B(N1482), .Y(N4040_1) );
  AND2X1 gate815 ( .A(N3691), .B(N4040_1), .Y(N4040) );
  AND2X1 gate816 ( .A(N3830), .B(N1583), .Y(N4041) );
  AND2X1 gate817 ( .A(N3831), .B(N1583), .Y(N4042) );
  AND2X1 gate818 ( .A(N3732), .B(N514), .Y(N4067) );
  AND2X1 gate819 ( .A(N514), .B(N3732), .Y(N4080) );
  AND2X1 gate820 ( .A(N3834), .B(N3668), .Y(N4088) );
  AND2X1 gate821 ( .A(N3835), .B(N3669), .Y(N4091) );
  AND2X1 gate822 ( .A(N3836), .B(N3670), .Y(N4094) );
  AND2X1 gate823 ( .A(N3837), .B(N3671), .Y(N4097) );
  AND2X1 gate824 ( .A(N3838), .B(N3676), .Y(N4100) );
  AND2X1 gate825 ( .A(N3839), .B(N3677), .Y(N4103) );
  AND2X1 gate826 ( .A(N3840), .B(N3678), .Y(N4106) );
  AND2X1 gate827 ( .A(N3841), .B(N3679), .Y(N4109) );
  AND2X1 gate828 ( .A(N3908), .B(N3703), .Y(N4144) );
  AND2X1 gate829 ( .A(N3909), .B(N3704), .Y(N4147) );
  BUFX2 gate830 ( .A(N3705), .Y(N4150) );
  AND2X1 gate831 ( .A(N3914), .B(N3711), .Y(N4153) );
  AND2X1 gate832 ( .A(N3915), .B(N3712), .Y(N4156) );
  AND2X1 gate833 ( .A(N3916), .B(N3713), .Y(N4159) );
  OR2X1 gate834 ( .A(N3758), .B(N3980), .Y(N4183) );
  OR2X1 gate835 ( .A(N3760), .B(N3981), .Y(N4184) );
  OR2X1 gate836_1 ( .A(N3761), .B(N3982), .Y(N4185_1) );
  OR2X1 gate836 ( .A(N446), .B(N4185_1), .Y(N4185) );
  OR2X1 gate837_1 ( .A(N3762), .B(N3983), .Y(N4186_1) );
  OR2X1 gate837 ( .A(N446), .B(N4186_1), .Y(N4186) );
  INVX1 gate838 ( .A(N3771), .Y(N4188) );
  INVX1 gate839 ( .A(N3775), .Y(N4191) );
  AND2X1 gate840_1 ( .A(N3775), .B(N3771), .Y(N4196_1) );
  AND2X1 gate840 ( .A(N3035), .B(N4196_1), .Y(N4196) );
  AND2X1 gate841_1 ( .A(N3987), .B(N3119), .Y(N4197_1) );
  AND2X1 gate841 ( .A(N3130), .B(N4197_1), .Y(N4197) );
  AND2X1 gate842 ( .A(N3920), .B(N3722), .Y(N4198) );
  INVX1 gate843 ( .A(N3816), .Y(N4199) );
  INVX1 gate844 ( .A(N3789), .Y(N4200) );
  INVX1 gate845 ( .A(N3793), .Y(N4203) );
  BUFX2 gate846 ( .A(N3797), .Y(N4206) );
  BUFX2 gate847 ( .A(N3797), .Y(N4209) );
  BUFX2 gate848 ( .A(N3732), .Y(N4212) );
  BUFX2 gate849 ( .A(N3732), .Y(N4215) );
  BUFX2 gate850 ( .A(N3732), .Y(N4219) );
  INVX1 gate851 ( .A(N3810), .Y(N4223) );
  INVX1 gate852 ( .A(N3813), .Y(N4224) );
  AND2X1 gate853 ( .A(N3918), .B(N3720), .Y(N4225) );
  AND2X1 gate854 ( .A(N3919), .B(N3721), .Y(N4228) );
  AND2X1 gate855 ( .A(N3991), .B(N3770), .Y(N4231) );
  AND2X1 gate856 ( .A(N3917), .B(N3719), .Y(N4234) );
  AND2X1 gate857 ( .A(N3989), .B(N3768), .Y(N4237) );
  AND2X1 gate858 ( .A(N3990), .B(N3769), .Y(N4240) );
  AND2X1 gate859 ( .A(N3988), .B(N3767), .Y(N4243) );
  AND2X1 gate860 ( .A(N3976), .B(N3746), .Y(N4246) );
  AND2X1 gate861 ( .A(N3977), .B(N3747), .Y(N4249) );
  AND2X1 gate862 ( .A(N3975), .B(N3745), .Y(N4252) );
  AND2X1 gate863 ( .A(N3978), .B(N3751), .Y(N4255) );
  AND2X1 gate864 ( .A(N3979), .B(N3752), .Y(N4258) );
  INVX1 gate865 ( .A(N3819), .Y(N4263) );
  NAND2X1 gate866 ( .A(N4024), .B(N3823), .Y(N4264) );
  INVX1 gate867 ( .A(N3824), .Y(N4267) );
  AND2X1 gate868 ( .A(N446), .B(N3893), .Y(N4268) );
  INVX1 gate869 ( .A(N3911), .Y(N4269) );
  INVX1 gate870 ( .A(N3984), .Y(N4270) );
  AND2X1 gate871 ( .A(N3893), .B(N446), .Y(N4271) );
  INVX1 gate872 ( .A(N4031), .Y(N4272) );
  OR2X1 gate873_1 ( .A(N4032), .B(N4033), .Y(N4273_1) );
  OR2X1 gate873_2 ( .A(N3614), .B(N3615), .Y(N4273_2) );
  OR2X1 gate873 ( .A(N4273_1), .B(N4273_2), .Y(N4273) );
  OR2X1 gate874_1 ( .A(N4034), .B(N4035), .Y(N4274_1) );
  OR2X1 gate874_2 ( .A(N3625), .B(N3626), .Y(N4274_2) );
  OR2X1 gate874 ( .A(N4274_1), .B(N4274_2), .Y(N4274) );
  INVX1 gate875 ( .A(N4036), .Y(N4275) );
  OR2X1 gate876_1 ( .A(N4037), .B(N4038), .Y(N4276_1) );
  OR2X1 gate876_2 ( .A(N3636), .B(N3637), .Y(N4276_2) );
  OR2X1 gate876 ( .A(N4276_1), .B(N4276_2), .Y(N4276) );
  OR2X1 gate877_1 ( .A(N4039), .B(N4040), .Y(N4277_1) );
  OR2X1 gate877_2 ( .A(N3639), .B(N3640), .Y(N4277_2) );
  OR2X1 gate877 ( .A(N4277_1), .B(N4277_2), .Y(N4277) );
  INVX1 gate878 ( .A(N4041), .Y(N4278) );
  INVX1 gate879 ( .A(N4042), .Y(N4279) );
  AND2X1 gate880 ( .A(N3887), .B(N457), .Y(N4280) );
  AND2X1 gate881 ( .A(N3881), .B(N468), .Y(N4284) );
  AND2X1 gate882 ( .A(N422), .B(N3873), .Y(N4290) );
  AND2X1 gate883 ( .A(N3867), .B(N435), .Y(N4297) );
  AND2X1 gate884 ( .A(N3861), .B(N389), .Y(N4298) );
  AND2X1 gate885 ( .A(N3855), .B(N400), .Y(N4301) );
  AND2X1 gate886 ( .A(N3849), .B(N411), .Y(N4305) );
  AND2X1 gate887 ( .A(N3842), .B(N374), .Y(N4310) );
  AND2X1 gate888 ( .A(N457), .B(N3887), .Y(N4316) );
  AND2X1 gate889 ( .A(N468), .B(N3881), .Y(N4320) );
  AND2X1 gate890 ( .A(N422), .B(N3873), .Y(N4325) );
  AND2X1 gate891 ( .A(N435), .B(N3867), .Y(N4331) );
  AND2X1 gate892 ( .A(N389), .B(N3861), .Y(N4332) );
  AND2X1 gate893 ( .A(N400), .B(N3855), .Y(N4336) );
  AND2X1 gate894 ( .A(N411), .B(N3849), .Y(N4342) );
  AND2X1 gate895 ( .A(N374), .B(N3842), .Y(N4349) );
  INVX1 gate896 ( .A(N3968), .Y(N4357) );
  INVX1 gate897 ( .A(N3962), .Y(N4364) );
  BUFX2 gate898 ( .A(N3962), .Y(N4375) );
  AND2X1 gate899 ( .A(N3956), .B(N479), .Y(N4379) );
  AND2X1 gate900 ( .A(N490), .B(N3948), .Y(N4385) );
  AND2X1 gate901 ( .A(N3942), .B(N503), .Y(N4392) );
  AND2X1 gate902 ( .A(N3933), .B(N523), .Y(N4396) );
  AND2X1 gate903 ( .A(N3927), .B(N534), .Y(N4400) );
  INVX1 gate904 ( .A(N3921), .Y(N4405) );
  BUFX2 gate905 ( .A(N3921), .Y(N4412) );
  INVX1 gate906 ( .A(N3968), .Y(N4418) );
  INVX1 gate907 ( .A(N3962), .Y(N4425) );
  BUFX2 gate908 ( .A(N3962), .Y(N4436) );
  AND2X1 gate909 ( .A(N479), .B(N3956), .Y(N4440) );
  AND2X1 gate910 ( .A(N490), .B(N3948), .Y(N4445) );
  AND2X1 gate911 ( .A(N503), .B(N3942), .Y(N4451) );
  AND2X1 gate912 ( .A(N523), .B(N3933), .Y(N4456) );
  AND2X1 gate913 ( .A(N534), .B(N3927), .Y(N4462) );
  BUFX2 gate914 ( .A(N3921), .Y(N4469) );
  INVX1 gate915 ( .A(N3921), .Y(N4477) );
  BUFX2 gate916 ( .A(N3968), .Y(N4512) );
  INVX1 gate917 ( .A(N4183), .Y(N4515) );
  INVX1 gate918 ( .A(N4184), .Y(N4516) );
  INVX1 gate919 ( .A(N4008), .Y(N4521) );
  INVX1 gate920 ( .A(N4011), .Y(N4523) );
  INVX1 gate921 ( .A(N4198), .Y(N4524) );
  INVX1 gate922 ( .A(N3984), .Y(N4532) );
  AND2X1 gate923_1 ( .A(N3911), .B(N3169), .Y(N4547_1) );
  AND2X1 gate923 ( .A(N3180), .B(N4547_1), .Y(N4547) );
  BUFX2 gate924 ( .A(N3893), .Y(N4548) );
  BUFX2 gate925 ( .A(N3887), .Y(N4551) );
  BUFX2 gate926 ( .A(N3881), .Y(N4554) );
  BUFX2 gate927 ( .A(N3873), .Y(N4557) );
  BUFX2 gate928 ( .A(N3867), .Y(N4560) );
  BUFX2 gate929 ( .A(N3861), .Y(N4563) );
  BUFX2 gate930 ( .A(N3855), .Y(N4566) );
  BUFX2 gate931 ( .A(N3849), .Y(N4569) );
  BUFX2 gate932 ( .A(N3842), .Y(N4572) );
  NOR2X1 gate933 ( .A(N422), .B(N3873), .Y(N4575) );
  BUFX2 gate934 ( .A(N3893), .Y(N4578) );
  BUFX2 gate935 ( .A(N3887), .Y(N4581) );
  BUFX2 gate936 ( .A(N3881), .Y(N4584) );
  BUFX2 gate937 ( .A(N3867), .Y(N4587) );
  BUFX2 gate938 ( .A(N3861), .Y(N4590) );
  BUFX2 gate939 ( .A(N3855), .Y(N4593) );
  BUFX2 gate940 ( .A(N3849), .Y(N4596) );
  BUFX2 gate941 ( .A(N3873), .Y(N4599) );
  BUFX2 gate942 ( .A(N3842), .Y(N4602) );
  NOR2X1 gate943 ( .A(N422), .B(N3873), .Y(N4605) );
  NOR2X1 gate944 ( .A(N374), .B(N3842), .Y(N4608) );
  BUFX2 gate945 ( .A(N3956), .Y(N4611) );
  BUFX2 gate946 ( .A(N3948), .Y(N4614) );
  BUFX2 gate947 ( .A(N3942), .Y(N4617) );
  BUFX2 gate948 ( .A(N3933), .Y(N4621) );
  BUFX2 gate949 ( .A(N3927), .Y(N4624) );
  NOR2X1 gate950 ( .A(N490), .B(N3948), .Y(N4627) );
  BUFX2 gate951 ( .A(N3956), .Y(N4630) );
  BUFX2 gate952 ( .A(N3942), .Y(N4633) );
  BUFX2 gate953 ( .A(N3933), .Y(N4637) );
  BUFX2 gate954 ( .A(N3927), .Y(N4640) );
  BUFX2 gate955 ( .A(N3948), .Y(N4643) );
  NOR2X1 gate956 ( .A(N490), .B(N3948), .Y(N4646) );
  BUFX2 gate957 ( .A(N3927), .Y(N4649) );
  BUFX2 gate958 ( .A(N3933), .Y(N4652) );
  BUFX2 gate959 ( .A(N3921), .Y(N4655) );
  BUFX2 gate960 ( .A(N3942), .Y(N4658) );
  BUFX2 gate961 ( .A(N3956), .Y(N4662) );
  BUFX2 gate962 ( .A(N3948), .Y(N4665) );
  BUFX2 gate963 ( .A(N3968), .Y(N4668) );
  BUFX2 gate964 ( .A(N3962), .Y(N4671) );
  BUFX2 gate965 ( .A(N3873), .Y(N4674) );
  BUFX2 gate966 ( .A(N3867), .Y(N4677) );
  BUFX2 gate967 ( .A(N3887), .Y(N4680) );
  BUFX2 gate968 ( .A(N3881), .Y(N4683) );
  BUFX2 gate969 ( .A(N3893), .Y(N4686) );
  BUFX2 gate970 ( .A(N3849), .Y(N4689) );
  BUFX2 gate971 ( .A(N3842), .Y(N4692) );
  BUFX2 gate972 ( .A(N3861), .Y(N4695) );
  BUFX2 gate973 ( .A(N3855), .Y(N4698) );
  NAND2X1 gate974 ( .A(N3813), .B(N4223), .Y(N4701) );
  NAND2X1 gate975 ( .A(N3810), .B(N4224), .Y(N4702) );
  INVX1 gate976 ( .A(N4021), .Y(N4720) );
  NAND2X1 gate977 ( .A(N4021), .B(N4263), .Y(N4721) );
  INVX1 gate978 ( .A(N4147), .Y(N4724) );
  INVX1 gate979 ( .A(N4144), .Y(N4725) );
  INVX1 gate980 ( .A(N4159), .Y(N4726) );
  INVX1 gate981 ( .A(N4156), .Y(N4727) );
  INVX1 gate982 ( .A(N4153), .Y(N4728) );
  INVX1 gate983 ( .A(N4097), .Y(N4729) );
  INVX1 gate984 ( .A(N4094), .Y(N4730) );
  INVX1 gate985 ( .A(N4091), .Y(N4731) );
  INVX1 gate986 ( .A(N4088), .Y(N4732) );
  INVX1 gate987 ( .A(N4109), .Y(N4733) );
  INVX1 gate988 ( .A(N4106), .Y(N4734) );
  INVX1 gate989 ( .A(N4103), .Y(N4735) );
  INVX1 gate990 ( .A(N4100), .Y(N4736) );
  AND2X1 gate991 ( .A(N4273), .B(N2877), .Y(N4737) );
  AND2X1 gate992 ( .A(N4274), .B(N2877), .Y(N4738) );
  AND2X1 gate993 ( .A(N4276), .B(N2877), .Y(N4739) );
  AND2X1 gate994 ( .A(N4277), .B(N2877), .Y(N4740) );
  AND2X1 gate995_1 ( .A(N4150), .B(N1758), .Y(N4741_1) );
  AND2X1 gate995 ( .A(N1755), .B(N4741_1), .Y(N4741) );
  INVX1 gate996 ( .A(N4212), .Y(N4855) );
  NAND2X1 gate997 ( .A(N4212), .B(N2712), .Y(N4856) );
  NAND2X1 gate998 ( .A(N4215), .B(N2718), .Y(N4908) );
  INVX1 gate999 ( .A(N4215), .Y(N4909) );
  AND2X1 gate1000 ( .A(N4515), .B(N4185), .Y(N4939) );
  AND2X1 gate1001 ( .A(N4516), .B(N4186), .Y(N4942) );
  INVX1 gate1002 ( .A(N4219), .Y(N4947) );
  AND2X1 gate1003_1 ( .A(N4188), .B(N3775), .Y(N4953_1) );
  AND2X1 gate1003 ( .A(N3779), .B(N4953_1), .Y(N4953) );
  AND2X1 gate1004_1 ( .A(N3771), .B(N4191), .Y(N4954_1) );
  AND2X1 gate1004 ( .A(N3780), .B(N4954_1), .Y(N4954) );
  AND2X1 gate1005_1 ( .A(N4191), .B(N4188), .Y(N4955_1) );
  AND2X1 gate1005 ( .A(N3038), .B(N4955_1), .Y(N4955) );
  AND2X1 gate1006_1 ( .A(N4109), .B(N3097), .Y(N4956_1) );
  AND2X1 gate1006 ( .A(N3108), .B(N4956_1), .Y(N4956) );
  AND2X1 gate1007_1 ( .A(N4106), .B(N3097), .Y(N4957_1) );
  AND2X1 gate1007 ( .A(N3108), .B(N4957_1), .Y(N4957) );
  AND2X1 gate1008_1 ( .A(N4103), .B(N3097), .Y(N4958_1) );
  AND2X1 gate1008 ( .A(N3108), .B(N4958_1), .Y(N4958) );
  AND2X1 gate1009_1 ( .A(N4100), .B(N3097), .Y(N4959_1) );
  AND2X1 gate1009 ( .A(N3108), .B(N4959_1), .Y(N4959) );
  AND2X1 gate1010_1 ( .A(N4159), .B(N3119), .Y(N4960_1) );
  AND2X1 gate1010 ( .A(N3130), .B(N4960_1), .Y(N4960) );
  AND2X1 gate1011_1 ( .A(N4156), .B(N3119), .Y(N4961_1) );
  AND2X1 gate1011 ( .A(N3130), .B(N4961_1), .Y(N4961) );
  INVX1 gate1012 ( .A(N4225), .Y(N4965) );
  INVX1 gate1013 ( .A(N4228), .Y(N4966) );
  INVX1 gate1014 ( .A(N4231), .Y(N4967) );
  INVX1 gate1015 ( .A(N4234), .Y(N4968) );
  INVX1 gate1016 ( .A(N4246), .Y(N4972) );
  INVX1 gate1017 ( .A(N4249), .Y(N4973) );
  INVX1 gate1018 ( .A(N4252), .Y(N4974) );
  NAND2X1 gate1019 ( .A(N4252), .B(N4199), .Y(N4975) );
  INVX1 gate1020 ( .A(N4206), .Y(N4976) );
  INVX1 gate1021 ( .A(N4209), .Y(N4977) );
  AND2X1 gate1022_1 ( .A(N3793), .B(N3789), .Y(N4978_1) );
  AND2X1 gate1022 ( .A(N4206), .B(N4978_1), .Y(N4978) );
  AND2X1 gate1023_1 ( .A(N4203), .B(N4200), .Y(N4979_1) );
  AND2X1 gate1023 ( .A(N4209), .B(N4979_1), .Y(N4979) );
  AND2X1 gate1024_1 ( .A(N4097), .B(N3147), .Y(N4980_1) );
  AND2X1 gate1024 ( .A(N3158), .B(N4980_1), .Y(N4980) );
  AND2X1 gate1025_1 ( .A(N4094), .B(N3147), .Y(N4981_1) );
  AND2X1 gate1025 ( .A(N3158), .B(N4981_1), .Y(N4981) );
  AND2X1 gate1026_1 ( .A(N4091), .B(N3147), .Y(N4982_1) );
  AND2X1 gate1026 ( .A(N3158), .B(N4982_1), .Y(N4982) );
  AND2X1 gate1027_1 ( .A(N4088), .B(N3147), .Y(N4983_1) );
  AND2X1 gate1027 ( .A(N3158), .B(N4983_1), .Y(N4983) );
  AND2X1 gate1028_1 ( .A(N4153), .B(N3169), .Y(N4984_1) );
  AND2X1 gate1028 ( .A(N3180), .B(N4984_1), .Y(N4984) );
  AND2X1 gate1029_1 ( .A(N4147), .B(N3169), .Y(N4985_1) );
  AND2X1 gate1029 ( .A(N3180), .B(N4985_1), .Y(N4985) );
  AND2X1 gate1030_1 ( .A(N4144), .B(N3169), .Y(N4986_1) );
  AND2X1 gate1030 ( .A(N3180), .B(N4986_1), .Y(N4986) );
  AND2X1 gate1031_1 ( .A(N4150), .B(N3169), .Y(N4987_1) );
  AND2X1 gate1031 ( .A(N3180), .B(N4987_1), .Y(N4987) );
  NAND2X1 gate1032 ( .A(N4701), .B(N4702), .Y(N5049) );
  INVX1 gate1033 ( .A(N4237), .Y(N5052) );
  INVX1 gate1034 ( .A(N4240), .Y(N5053) );
  INVX1 gate1035 ( .A(N4243), .Y(N5054) );
  INVX1 gate1036 ( .A(N4255), .Y(N5055) );
  INVX1 gate1037 ( .A(N4258), .Y(N5056) );
  NAND2X1 gate1038 ( .A(N3819), .B(N4720), .Y(N5057) );
  INVX1 gate1039 ( .A(N4264), .Y(N5058) );
  NAND2X1 gate1040 ( .A(N4264), .B(N4267), .Y(N5059) );
  AND2X1 gate1041_1 ( .A(N4724), .B(N4725), .Y(N5060_1) );
  AND2X1 gate1041_2 ( .A(N4269), .B(N4027), .Y(N5060_2) );
  AND2X1 gate1041 ( .A(N5060_1), .B(N5060_2), .Y(N5060) );
  AND2X1 gate1042_1 ( .A(N4726), .B(N4727), .Y(N5061_1) );
  AND2X1 gate1042_2 ( .A(N3827), .B(N4728), .Y(N5061_2) );
  AND2X1 gate1042 ( .A(N5061_1), .B(N5061_2), .Y(N5061) );
  AND2X1 gate1043_1 ( .A(N4729), .B(N4730), .Y(N5062_1) );
  AND2X1 gate1043_2 ( .A(N4731), .B(N4732), .Y(N5062_2) );
  AND2X1 gate1043 ( .A(N5062_1), .B(N5062_2), .Y(N5062) );
  AND2X1 gate1044_1 ( .A(N4733), .B(N4734), .Y(N5063_1) );
  AND2X1 gate1044_2 ( .A(N4735), .B(N4736), .Y(N5063_2) );
  AND2X1 gate1044 ( .A(N5063_1), .B(N5063_2), .Y(N5063) );
  AND2X1 gate1045 ( .A(N4357), .B(N4375), .Y(N5065) );
  AND2X1 gate1046_1 ( .A(N4364), .B(N4357), .Y(N5066_1) );
  AND2X1 gate1046 ( .A(N4379), .B(N5066_1), .Y(N5066) );
  AND2X1 gate1047 ( .A(N4418), .B(N4436), .Y(N5067) );
  AND2X1 gate1048_1 ( .A(N4425), .B(N4418), .Y(N5068_1) );
  AND2X1 gate1048 ( .A(N4440), .B(N5068_1), .Y(N5068) );
  INVX1 gate1049 ( .A(N4548), .Y(N5069) );
  NAND2X1 gate1050 ( .A(N4548), .B(N2628), .Y(N5070) );
  INVX1 gate1051 ( .A(N4551), .Y(N5071) );
  NAND2X1 gate1052 ( .A(N4551), .B(N2629), .Y(N5072) );
  INVX1 gate1053 ( .A(N4554), .Y(N5073) );
  NAND2X1 gate1054 ( .A(N4554), .B(N2630), .Y(N5074) );
  INVX1 gate1055 ( .A(N4557), .Y(N5075) );
  NAND2X1 gate1056 ( .A(N4557), .B(N2631), .Y(N5076) );
  INVX1 gate1057 ( .A(N4560), .Y(N5077) );
  NAND2X1 gate1058 ( .A(N4560), .B(N2632), .Y(N5078) );
  INVX1 gate1059 ( .A(N4563), .Y(N5079) );
  NAND2X1 gate1060 ( .A(N4563), .B(N2633), .Y(N5080) );
  INVX1 gate1061 ( .A(N4566), .Y(N5081) );
  NAND2X1 gate1062 ( .A(N4566), .B(N2634), .Y(N5082) );
  INVX1 gate1063 ( .A(N4569), .Y(N5083) );
  NAND2X1 gate1064 ( .A(N4569), .B(N2635), .Y(N5084) );
  INVX1 gate1065 ( .A(N4572), .Y(N5085) );
  NAND2X1 gate1066 ( .A(N4572), .B(N2636), .Y(N5086) );
  INVX1 gate1067 ( .A(N4575), .Y(N5087) );
  NAND2X1 gate1068 ( .A(N4578), .B(N2638), .Y(N5088) );
  INVX1 gate1069 ( .A(N4578), .Y(N5089) );
  NAND2X1 gate1070 ( .A(N4581), .B(N2639), .Y(N5090) );
  INVX1 gate1071 ( .A(N4581), .Y(N5091) );
  NAND2X1 gate1072 ( .A(N4584), .B(N2640), .Y(N5092) );
  INVX1 gate1073 ( .A(N4584), .Y(N5093) );
  NAND2X1 gate1074 ( .A(N4587), .B(N2641), .Y(N5094) );
  INVX1 gate1075 ( .A(N4587), .Y(N5095) );
  NAND2X1 gate1076 ( .A(N4590), .B(N2642), .Y(N5096) );
  INVX1 gate1077 ( .A(N4590), .Y(N5097) );
  NAND2X1 gate1078 ( .A(N4593), .B(N2643), .Y(N5098) );
  INVX1 gate1079 ( .A(N4593), .Y(N5099) );
  NAND2X1 gate1080 ( .A(N4596), .B(N2644), .Y(N5100) );
  INVX1 gate1081 ( .A(N4596), .Y(N5101) );
  NAND2X1 gate1082 ( .A(N4599), .B(N2645), .Y(N5102) );
  INVX1 gate1083 ( .A(N4599), .Y(N5103) );
  NAND2X1 gate1084 ( .A(N4602), .B(N2646), .Y(N5104) );
  INVX1 gate1085 ( .A(N4602), .Y(N5105) );
  INVX1 gate1086 ( .A(N4611), .Y(N5106) );
  NAND2X1 gate1087 ( .A(N4611), .B(N2709), .Y(N5107) );
  INVX1 gate1088 ( .A(N4614), .Y(N5108) );
  NAND2X1 gate1089 ( .A(N4614), .B(N2710), .Y(N5109) );
  INVX1 gate1090 ( .A(N4617), .Y(N5110) );
  NAND2X1 gate1091 ( .A(N4617), .B(N2711), .Y(N5111) );
  NAND2X1 gate1092 ( .A(N1890), .B(N4855), .Y(N5112) );
  INVX1 gate1093 ( .A(N4621), .Y(N5113) );
  NAND2X1 gate1094 ( .A(N4621), .B(N2713), .Y(N5114) );
  INVX1 gate1095 ( .A(N4624), .Y(N5115) );
  NAND2X1 gate1096 ( .A(N4624), .B(N2714), .Y(N5116) );
  AND2X1 gate1097 ( .A(N4364), .B(N4379), .Y(N5117) );
  AND2X1 gate1098 ( .A(N4364), .B(N4379), .Y(N5118) );
  AND2X1 gate1099 ( .A(N54), .B(N4405), .Y(N5119) );
  INVX1 gate1100 ( .A(N4627), .Y(N5120) );
  NAND2X1 gate1101 ( .A(N4630), .B(N2716), .Y(N5121) );
  INVX1 gate1102 ( .A(N4630), .Y(N5122) );
  NAND2X1 gate1103 ( .A(N4633), .B(N2717), .Y(N5123) );
  INVX1 gate1104 ( .A(N4633), .Y(N5124) );
  NAND2X1 gate1105 ( .A(N1908), .B(N4909), .Y(N5125) );
  NAND2X1 gate1106 ( .A(N4637), .B(N2719), .Y(N5126) );
  INVX1 gate1107 ( .A(N4637), .Y(N5127) );
  NAND2X1 gate1108 ( .A(N4640), .B(N2720), .Y(N5128) );
  INVX1 gate1109 ( .A(N4640), .Y(N5129) );
  NAND2X1 gate1110 ( .A(N4643), .B(N2721), .Y(N5130) );
  INVX1 gate1111 ( .A(N4643), .Y(N5131) );
  AND2X1 gate1112 ( .A(N4425), .B(N4440), .Y(N5132) );
  AND2X1 gate1113 ( .A(N4425), .B(N4440), .Y(N5133) );
  INVX1 gate1114 ( .A(N4649), .Y(N5135) );
  INVX1 gate1115 ( .A(N4652), .Y(N5136) );
  NAND2X1 gate1116 ( .A(N4655), .B(N4521), .Y(N5137) );
  INVX1 gate1117 ( .A(N4655), .Y(N5138) );
  INVX1 gate1118 ( .A(N4658), .Y(N5139) );
  NAND2X1 gate1119 ( .A(N4658), .B(N4947), .Y(N5140) );
  INVX1 gate1120 ( .A(N4674), .Y(N5141) );
  INVX1 gate1121 ( .A(N4677), .Y(N5142) );
  INVX1 gate1122 ( .A(N4680), .Y(N5143) );
  INVX1 gate1123 ( .A(N4683), .Y(N5144) );
  NAND2X1 gate1124 ( .A(N4686), .B(N4523), .Y(N5145) );
  INVX1 gate1125 ( .A(N4686), .Y(N5146) );
  NOR2X1 gate1126 ( .A(N4953), .B(N4196), .Y(N5147) );
  NOR2X1 gate1127 ( .A(N4954), .B(N4955), .Y(N5148) );
  INVX1 gate1128 ( .A(N4524), .Y(N5150) );
  NAND2X1 gate1129 ( .A(N4228), .B(N4965), .Y(N5153) );
  NAND2X1 gate1130 ( .A(N4225), .B(N4966), .Y(N5154) );
  NAND2X1 gate1131 ( .A(N4234), .B(N4967), .Y(N5155) );
  NAND2X1 gate1132 ( .A(N4231), .B(N4968), .Y(N5156) );
  INVX1 gate1133 ( .A(N4532), .Y(N5157) );
  NAND2X1 gate1134 ( .A(N4249), .B(N4972), .Y(N5160) );
  NAND2X1 gate1135 ( .A(N4246), .B(N4973), .Y(N5161) );
  NAND2X1 gate1136 ( .A(N3816), .B(N4974), .Y(N5162) );
  AND2X1 gate1137_1 ( .A(N4200), .B(N3793), .Y(N5163_1) );
  AND2X1 gate1137 ( .A(N4976), .B(N5163_1), .Y(N5163) );
  AND2X1 gate1138_1 ( .A(N3789), .B(N4203), .Y(N5164_1) );
  AND2X1 gate1138 ( .A(N4977), .B(N5164_1), .Y(N5164) );
  AND2X1 gate1139_1 ( .A(N4942), .B(N3147), .Y(N5165_1) );
  AND2X1 gate1139 ( .A(N3158), .B(N5165_1), .Y(N5165) );
  INVX1 gate1140 ( .A(N4512), .Y(N5166) );
  BUFX2 gate1141 ( .A(N4290), .Y(N5169) );
  INVX1 gate1142 ( .A(N4605), .Y(N5172) );
  BUFX2 gate1143 ( .A(N4325), .Y(N5173) );
  INVX1 gate1144 ( .A(N4608), .Y(N5176) );
  BUFX2 gate1145 ( .A(N4349), .Y(N5177) );
  BUFX2 gate1146 ( .A(N4405), .Y(N5180) );
  BUFX2 gate1147 ( .A(N4357), .Y(N5183) );
  BUFX2 gate1148 ( .A(N4357), .Y(N5186) );
  BUFX2 gate1149 ( .A(N4364), .Y(N5189) );
  BUFX2 gate1150 ( .A(N4364), .Y(N5192) );
  BUFX2 gate1151 ( .A(N4385), .Y(N5195) );
  INVX1 gate1152 ( .A(N4646), .Y(N5198) );
  BUFX2 gate1153 ( .A(N4418), .Y(N5199) );
  BUFX2 gate1154 ( .A(N4425), .Y(N5202) );
  BUFX2 gate1155 ( .A(N4445), .Y(N5205) );
  BUFX2 gate1156 ( .A(N4418), .Y(N5208) );
  BUFX2 gate1157 ( .A(N4425), .Y(N5211) );
  BUFX2 gate1158 ( .A(N4477), .Y(N5214) );
  BUFX2 gate1159 ( .A(N4469), .Y(N5217) );
  BUFX2 gate1160 ( .A(N4477), .Y(N5220) );
  INVX1 gate1161 ( .A(N4662), .Y(N5223) );
  INVX1 gate1162 ( .A(N4665), .Y(N5224) );
  INVX1 gate1163 ( .A(N4668), .Y(N5225) );
  INVX1 gate1164 ( .A(N4671), .Y(N5226) );
  INVX1 gate1165 ( .A(N4689), .Y(N5227) );
  INVX1 gate1166 ( .A(N4692), .Y(N5228) );
  INVX1 gate1167 ( .A(N4695), .Y(N5229) );
  INVX1 gate1168 ( .A(N4698), .Y(N5230) );
  NAND2X1 gate1169 ( .A(N4240), .B(N5052), .Y(N5232) );
  NAND2X1 gate1170 ( .A(N4237), .B(N5053), .Y(N5233) );
  NAND2X1 gate1171 ( .A(N4258), .B(N5055), .Y(N5234) );
  NAND2X1 gate1172 ( .A(N4255), .B(N5056), .Y(N5235) );
  NAND2X1 gate1173 ( .A(N4721), .B(N5057), .Y(N5236) );
  NAND2X1 gate1174 ( .A(N3824), .B(N5058), .Y(N5239) );
  AND2X1 gate1175_1 ( .A(N5060), .B(N5061), .Y(N5240_1) );
  AND2X1 gate1175 ( .A(N4270), .B(N5240_1), .Y(N5240) );
  INVX1 gate1176 ( .A(N4939), .Y(N5241) );
  NAND2X1 gate1177 ( .A(N1824), .B(N5069), .Y(N5242) );
  NAND2X1 gate1178 ( .A(N1827), .B(N5071), .Y(N5243) );
  NAND2X1 gate1179 ( .A(N1830), .B(N5073), .Y(N5244) );
  NAND2X1 gate1180 ( .A(N1833), .B(N5075), .Y(N5245) );
  NAND2X1 gate1181 ( .A(N1836), .B(N5077), .Y(N5246) );
  NAND2X1 gate1182 ( .A(N1839), .B(N5079), .Y(N5247) );
  NAND2X1 gate1183 ( .A(N1842), .B(N5081), .Y(N5248) );
  NAND2X1 gate1184 ( .A(N1845), .B(N5083), .Y(N5249) );
  NAND2X1 gate1185 ( .A(N1848), .B(N5085), .Y(N5250) );
  NAND2X1 gate1186 ( .A(N1854), .B(N5089), .Y(N5252) );
  NAND2X1 gate1187 ( .A(N1857), .B(N5091), .Y(N5253) );
  NAND2X1 gate1188 ( .A(N1860), .B(N5093), .Y(N5254) );
  NAND2X1 gate1189 ( .A(N1863), .B(N5095), .Y(N5255) );
  NAND2X1 gate1190 ( .A(N1866), .B(N5097), .Y(N5256) );
  NAND2X1 gate1191 ( .A(N1869), .B(N5099), .Y(N5257) );
  NAND2X1 gate1192 ( .A(N1872), .B(N5101), .Y(N5258) );
  NAND2X1 gate1193 ( .A(N1875), .B(N5103), .Y(N5259) );
  NAND2X1 gate1194 ( .A(N1878), .B(N5105), .Y(N5260) );
  NAND2X1 gate1195 ( .A(N1881), .B(N5106), .Y(N5261) );
  NAND2X1 gate1196 ( .A(N1884), .B(N5108), .Y(N5262) );
  NAND2X1 gate1197 ( .A(N1887), .B(N5110), .Y(N5263) );
  NAND2X1 gate1198 ( .A(N5112), .B(N4856), .Y(N5264) );
  NAND2X1 gate1199 ( .A(N1893), .B(N5113), .Y(N5274) );
  NAND2X1 gate1200 ( .A(N1896), .B(N5115), .Y(N5275) );
  NAND2X1 gate1201 ( .A(N1902), .B(N5122), .Y(N5282) );
  NAND2X1 gate1202 ( .A(N1905), .B(N5124), .Y(N5283) );
  NAND2X1 gate1203 ( .A(N4908), .B(N5125), .Y(N5284) );
  NAND2X1 gate1204 ( .A(N1911), .B(N5127), .Y(N5298) );
  NAND2X1 gate1205 ( .A(N1914), .B(N5129), .Y(N5299) );
  NAND2X1 gate1206 ( .A(N1917), .B(N5131), .Y(N5300) );
  NAND2X1 gate1207 ( .A(N4652), .B(N5135), .Y(N5303) );
  NAND2X1 gate1208 ( .A(N4649), .B(N5136), .Y(N5304) );
  NAND2X1 gate1209 ( .A(N4008), .B(N5138), .Y(N5305) );
  NAND2X1 gate1210 ( .A(N4219), .B(N5139), .Y(N5306) );
  NAND2X1 gate1211 ( .A(N4677), .B(N5141), .Y(N5307) );
  NAND2X1 gate1212 ( .A(N4674), .B(N5142), .Y(N5308) );
  NAND2X1 gate1213 ( .A(N4683), .B(N5143), .Y(N5309) );
  NAND2X1 gate1214 ( .A(N4680), .B(N5144), .Y(N5310) );
  NAND2X1 gate1215 ( .A(N4011), .B(N5146), .Y(N5311) );
  INVX1 gate1216 ( .A(N5049), .Y(N5312) );
  NAND2X1 gate1217 ( .A(N5153), .B(N5154), .Y(N5315) );
  NAND2X1 gate1218 ( .A(N5155), .B(N5156), .Y(N5319) );
  NAND2X1 gate1219 ( .A(N5160), .B(N5161), .Y(N5324) );
  NAND2X1 gate1220 ( .A(N5162), .B(N4975), .Y(N5328) );
  NOR2X1 gate1221 ( .A(N5163), .B(N4978), .Y(N5331) );
  NOR2X1 gate1222 ( .A(N5164), .B(N4979), .Y(N5332) );
  OR2X1 gate1223 ( .A(N4412), .B(N5119), .Y(N5346) );
  NAND2X1 gate1224 ( .A(N4665), .B(N5223), .Y(N5363) );
  NAND2X1 gate1225 ( .A(N4662), .B(N5224), .Y(N5364) );
  NAND2X1 gate1226 ( .A(N4671), .B(N5225), .Y(N5365) );
  NAND2X1 gate1227 ( .A(N4668), .B(N5226), .Y(N5366) );
  NAND2X1 gate1228 ( .A(N4692), .B(N5227), .Y(N5367) );
  NAND2X1 gate1229 ( .A(N4689), .B(N5228), .Y(N5368) );
  NAND2X1 gate1230 ( .A(N4698), .B(N5229), .Y(N5369) );
  NAND2X1 gate1231 ( .A(N4695), .B(N5230), .Y(N5370) );
  NAND2X1 gate1232 ( .A(N5148), .B(N5147), .Y(N5371) );
  BUFX2 gate1233 ( .A(N4939), .Y(N5374) );
  NAND2X1 gate1234 ( .A(N5232), .B(N5233), .Y(N5377) );
  NAND2X1 gate1235 ( .A(N5234), .B(N5235), .Y(N5382) );
  NAND2X1 gate1236 ( .A(N5239), .B(N5059), .Y(N5385) );
  AND2X1 gate1237_1 ( .A(N5062), .B(N5063), .Y(N5388_1) );
  AND2X1 gate1237 ( .A(N5241), .B(N5388_1), .Y(N5388) );
  NAND2X1 gate1238 ( .A(N5242), .B(N5070), .Y(N5389) );
  NAND2X1 gate1239 ( .A(N5243), .B(N5072), .Y(N5396) );
  NAND2X1 gate1240 ( .A(N5244), .B(N5074), .Y(N5407) );
  NAND2X1 gate1241 ( .A(N5245), .B(N5076), .Y(N5418) );
  NAND2X1 gate1242 ( .A(N5246), .B(N5078), .Y(N5424) );
  NAND2X1 gate1243 ( .A(N5247), .B(N5080), .Y(N5431) );
  NAND2X1 gate1244 ( .A(N5248), .B(N5082), .Y(N5441) );
  NAND2X1 gate1245 ( .A(N5249), .B(N5084), .Y(N5452) );
  NAND2X1 gate1246 ( .A(N5250), .B(N5086), .Y(N5462) );
  INVX1 gate1247 ( .A(N5169), .Y(N5469) );
  NAND2X1 gate1248 ( .A(N5088), .B(N5252), .Y(N5470) );
  NAND2X1 gate1249 ( .A(N5090), .B(N5253), .Y(N5477) );
  NAND2X1 gate1250 ( .A(N5092), .B(N5254), .Y(N5488) );
  NAND2X1 gate1251 ( .A(N5094), .B(N5255), .Y(N5498) );
  NAND2X1 gate1252 ( .A(N5096), .B(N5256), .Y(N5506) );
  NAND2X1 gate1253 ( .A(N5098), .B(N5257), .Y(N5520) );
  NAND2X1 gate1254 ( .A(N5100), .B(N5258), .Y(N5536) );
  NAND2X1 gate1255 ( .A(N5102), .B(N5259), .Y(N5549) );
  NAND2X1 gate1256 ( .A(N5104), .B(N5260), .Y(N5555) );
  NAND2X1 gate1257 ( .A(N5261), .B(N5107), .Y(N5562) );
  NAND2X1 gate1258 ( .A(N5262), .B(N5109), .Y(N5573) );
  NAND2X1 gate1259 ( .A(N5263), .B(N5111), .Y(N5579) );
  NAND2X1 gate1260 ( .A(N5274), .B(N5114), .Y(N5595) );
  NAND2X1 gate1261 ( .A(N5275), .B(N5116), .Y(N5606) );
  NAND2X1 gate1262 ( .A(N5180), .B(N2715), .Y(N5616) );
  INVX1 gate1263 ( .A(N5180), .Y(N5617) );
  INVX1 gate1264 ( .A(N5183), .Y(N5618) );
  INVX1 gate1265 ( .A(N5186), .Y(N5619) );
  INVX1 gate1266 ( .A(N5189), .Y(N5620) );
  INVX1 gate1267 ( .A(N5192), .Y(N5621) );
  INVX1 gate1268 ( .A(N5195), .Y(N5622) );
  NAND2X1 gate1269 ( .A(N5121), .B(N5282), .Y(N5624) );
  NAND2X1 gate1270 ( .A(N5123), .B(N5283), .Y(N5634) );
  NAND2X1 gate1271 ( .A(N5126), .B(N5298), .Y(N5655) );
  NAND2X1 gate1272 ( .A(N5128), .B(N5299), .Y(N5671) );
  NAND2X1 gate1273 ( .A(N5130), .B(N5300), .Y(N5684) );
  INVX1 gate1274 ( .A(N5202), .Y(N5690) );
  INVX1 gate1275 ( .A(N5211), .Y(N5691) );
  NAND2X1 gate1276 ( .A(N5303), .B(N5304), .Y(N5692) );
  NAND2X1 gate1277 ( .A(N5137), .B(N5305), .Y(N5696) );
  NAND2X1 gate1278 ( .A(N5306), .B(N5140), .Y(N5700) );
  NAND2X1 gate1279 ( .A(N5307), .B(N5308), .Y(N5703) );
  NAND2X1 gate1280 ( .A(N5309), .B(N5310), .Y(N5707) );
  NAND2X1 gate1281 ( .A(N5145), .B(N5311), .Y(N5711) );
  AND2X1 gate1282 ( .A(N5166), .B(N4512), .Y(N5726) );
  INVX1 gate1283 ( .A(N5173), .Y(N5727) );
  INVX1 gate1284 ( .A(N5177), .Y(N5728) );
  INVX1 gate1285 ( .A(N5199), .Y(N5730) );
  INVX1 gate1286 ( .A(N5205), .Y(N5731) );
  INVX1 gate1287 ( .A(N5208), .Y(N5732) );
  INVX1 gate1288 ( .A(N5214), .Y(N5733) );
  INVX1 gate1289 ( .A(N5217), .Y(N5734) );
  INVX1 gate1290 ( .A(N5220), .Y(N5735) );
  NAND2X1 gate1291 ( .A(N5365), .B(N5366), .Y(N5736) );
  NAND2X1 gate1292 ( .A(N5363), .B(N5364), .Y(N5739) );
  NAND2X1 gate1293 ( .A(N5369), .B(N5370), .Y(N5742) );
  NAND2X1 gate1294 ( .A(N5367), .B(N5368), .Y(N5745) );
  INVX1 gate1295 ( .A(N5236), .Y(N5755) );
  NAND2X1 gate1296 ( .A(N5332), .B(N5331), .Y(N5756) );
  AND2X1 gate1297 ( .A(N5264), .B(N4396), .Y(N5954) );
  NAND2X1 gate1298 ( .A(N1899), .B(N5617), .Y(N5955) );
  INVX1 gate1299 ( .A(N5346), .Y(N5956) );
  AND2X1 gate1300 ( .A(N5284), .B(N4456), .Y(N6005) );
  AND2X1 gate1301 ( .A(N5284), .B(N4456), .Y(N6006) );
  INVX1 gate1302 ( .A(N5371), .Y(N6023) );
  NAND2X1 gate1303 ( .A(N5371), .B(N5312), .Y(N6024) );
  INVX1 gate1304 ( .A(N5315), .Y(N6025) );
  INVX1 gate1305 ( .A(N5324), .Y(N6028) );
  BUFX2 gate1306 ( .A(N5319), .Y(N6031) );
  BUFX2 gate1307 ( .A(N5319), .Y(N6034) );
  BUFX2 gate1308 ( .A(N5328), .Y(N6037) );
  BUFX2 gate1309 ( .A(N5328), .Y(N6040) );
  INVX1 gate1310 ( .A(N5385), .Y(N6044) );
  OR2X1 gate1311 ( .A(N5166), .B(N5726), .Y(N6045) );
  BUFX2 gate1312 ( .A(N5264), .Y(N6048) );
  BUFX2 gate1313 ( .A(N5284), .Y(N6051) );
  BUFX2 gate1314 ( .A(N5284), .Y(N6054) );
  INVX1 gate1315 ( .A(N5374), .Y(N6065) );
  NAND2X1 gate1316 ( .A(N5374), .B(N5054), .Y(N6066) );
  INVX1 gate1317 ( .A(N5377), .Y(N6067) );
  INVX1 gate1318 ( .A(N5382), .Y(N6068) );
  NAND2X1 gate1319 ( .A(N5382), .B(N5755), .Y(N6069) );
  AND2X1 gate1320 ( .A(N5470), .B(N4316), .Y(N6071) );
  AND2X1 gate1321_1 ( .A(N5477), .B(N5470), .Y(N6072_1) );
  AND2X1 gate1321 ( .A(N4320), .B(N6072_1), .Y(N6072) );
  AND2X1 gate1322_1 ( .A(N5488), .B(N5470), .Y(N6073_1) );
  AND2X1 gate1322_2 ( .A(N4325), .B(N5477), .Y(N6073_2) );
  AND2X1 gate1322 ( .A(N6073_1), .B(N6073_2), .Y(N6073) );
  AND2X1 gate1323_1 ( .A(N5562), .B(N4357), .Y(N6074_1) );
  AND2X1 gate1323_2 ( .A(N4385), .B(N4364), .Y(N6074_2) );
  AND2X1 gate1323 ( .A(N6074_1), .B(N6074_2), .Y(N6074) );
  AND2X1 gate1324 ( .A(N5389), .B(N4280), .Y(N6075) );
  AND2X1 gate1325_1 ( .A(N5396), .B(N5389), .Y(N6076_1) );
  AND2X1 gate1325 ( .A(N4284), .B(N6076_1), .Y(N6076) );
  AND2X1 gate1326_1 ( .A(N5407), .B(N5389), .Y(N6077_1) );
  AND2X1 gate1326_2 ( .A(N4290), .B(N5396), .Y(N6077_2) );
  AND2X1 gate1326 ( .A(N6077_1), .B(N6077_2), .Y(N6077) );
  AND2X1 gate1327_1 ( .A(N5624), .B(N4418), .Y(N6078_1) );
  AND2X1 gate1327_2 ( .A(N4445), .B(N4425), .Y(N6078_2) );
  AND2X1 gate1327 ( .A(N6078_1), .B(N6078_2), .Y(N6078) );
  INVX1 gate1328 ( .A(N5418), .Y(N6079) );
  AND2X1 gate1329_1 ( .A(N5396), .B(N5418), .Y(N6080_1) );
  AND2X1 gate1329_2 ( .A(N5407), .B(N5389), .Y(N6080_2) );
  AND2X1 gate1329 ( .A(N6080_1), .B(N6080_2), .Y(N6080) );
  AND2X1 gate1330 ( .A(N5396), .B(N4284), .Y(N6083) );
  AND2X1 gate1331_1 ( .A(N5407), .B(N4290), .Y(N6084_1) );
  AND2X1 gate1331 ( .A(N5396), .B(N6084_1), .Y(N6084) );
  AND2X1 gate1332_1 ( .A(N5418), .B(N5407), .Y(N6085_1) );
  AND2X1 gate1332 ( .A(N5396), .B(N6085_1), .Y(N6085) );
  AND2X1 gate1333 ( .A(N5396), .B(N4284), .Y(N6086) );
  AND2X1 gate1334_1 ( .A(N4290), .B(N5407), .Y(N6087_1) );
  AND2X1 gate1334 ( .A(N5396), .B(N6087_1), .Y(N6087) );
  AND2X1 gate1335 ( .A(N5407), .B(N4290), .Y(N6088) );
  AND2X1 gate1336 ( .A(N5418), .B(N5407), .Y(N6089) );
  AND2X1 gate1337 ( .A(N5407), .B(N4290), .Y(N6090) );
  AND2X1 gate1338_1 ( .A(N5431), .B(N5462), .Y(N6091_1) );
  AND2X1 gate1338_2 ( .A(N5441), .B(N5424), .Y(N6091_2) );
  AND2X1 gate1338_3 ( .A(N5452), .B(N6091_1), .Y(N6091_3) );
  AND2X1 gate1338 ( .A(N6091_2), .B(N6091_3), .Y(N6091) );
  AND2X1 gate1339 ( .A(N5424), .B(N4298), .Y(N6094) );
  AND2X1 gate1340_1 ( .A(N5431), .B(N5424), .Y(N6095_1) );
  AND2X1 gate1340 ( .A(N4301), .B(N6095_1), .Y(N6095) );
  AND2X1 gate1341_1 ( .A(N5441), .B(N5424), .Y(N6096_1) );
  AND2X1 gate1341_2 ( .A(N4305), .B(N5431), .Y(N6096_2) );
  AND2X1 gate1341 ( .A(N6096_1), .B(N6096_2), .Y(N6096) );
  AND2X1 gate1342_1 ( .A(N5452), .B(N5441), .Y(N6097_1) );
  AND2X1 gate1342_2 ( .A(N5424), .B(N4310), .Y(N6097_2) );
  AND2X1 gate1342_3 ( .A(N5431), .B(N6097_1), .Y(N6097_3) );
  AND2X1 gate1342 ( .A(N6097_2), .B(N6097_3), .Y(N6097) );
  AND2X1 gate1343 ( .A(N5431), .B(N4301), .Y(N6098) );
  AND2X1 gate1344_1 ( .A(N5441), .B(N4305), .Y(N6099_1) );
  AND2X1 gate1344 ( .A(N5431), .B(N6099_1), .Y(N6099) );
  AND2X1 gate1345_1 ( .A(N5452), .B(N5441), .Y(N6100_1) );
  AND2X1 gate1345_2 ( .A(N4310), .B(N5431), .Y(N6100_2) );
  AND2X1 gate1345 ( .A(N6100_1), .B(N6100_2), .Y(N6100) );
  AND2X1 gate1346_1 ( .A(N4), .B(N5462), .Y(N6101_1) );
  AND2X1 gate1346_2 ( .A(N5441), .B(N5452), .Y(N6101_2) );
  AND2X1 gate1346_3 ( .A(N5431), .B(N6101_1), .Y(N6101_3) );
  AND2X1 gate1346 ( .A(N6101_2), .B(N6101_3), .Y(N6101) );
  AND2X1 gate1347 ( .A(N4305), .B(N5441), .Y(N6102) );
  AND2X1 gate1348_1 ( .A(N5452), .B(N5441), .Y(N6103_1) );
  AND2X1 gate1348 ( .A(N4310), .B(N6103_1), .Y(N6103) );
  AND2X1 gate1349_1 ( .A(N4), .B(N5462), .Y(N6104_1) );
  AND2X1 gate1349_2 ( .A(N5441), .B(N5452), .Y(N6104_2) );
  AND2X1 gate1349 ( .A(N6104_1), .B(N6104_2), .Y(N6104) );
  AND2X1 gate1350 ( .A(N5452), .B(N4310), .Y(N6105) );
  AND2X1 gate1351_1 ( .A(N4), .B(N5462), .Y(N6106_1) );
  AND2X1 gate1351 ( .A(N5452), .B(N6106_1), .Y(N6106) );
  AND2X1 gate1352 ( .A(N4), .B(N5462), .Y(N6107) );
  AND2X1 gate1353_1 ( .A(N5549), .B(N5488), .Y(N6108_1) );
  AND2X1 gate1353_2 ( .A(N5477), .B(N5470), .Y(N6108_2) );
  AND2X1 gate1353 ( .A(N6108_1), .B(N6108_2), .Y(N6108) );
  AND2X1 gate1354 ( .A(N5477), .B(N4320), .Y(N6111) );
  AND2X1 gate1355_1 ( .A(N5488), .B(N4325), .Y(N6112_1) );
  AND2X1 gate1355 ( .A(N5477), .B(N6112_1), .Y(N6112) );
  AND2X1 gate1356_1 ( .A(N5549), .B(N5488), .Y(N6113_1) );
  AND2X1 gate1356 ( .A(N5477), .B(N6113_1), .Y(N6113) );
  AND2X1 gate1357 ( .A(N5477), .B(N4320), .Y(N6114) );
  AND2X1 gate1358_1 ( .A(N5488), .B(N4325), .Y(N6115_1) );
  AND2X1 gate1358 ( .A(N5477), .B(N6115_1), .Y(N6115) );
  AND2X1 gate1359 ( .A(N5488), .B(N4325), .Y(N6116) );
  AND2X1 gate1360_1 ( .A(N5555), .B(N5536), .Y(N6117_1) );
  AND2X1 gate1360_2 ( .A(N5520), .B(N5506), .Y(N6117_2) );
  AND2X1 gate1360_3 ( .A(N5498), .B(N6117_1), .Y(N6117_3) );
  AND2X1 gate1360 ( .A(N6117_2), .B(N6117_3), .Y(N6117) );
  AND2X1 gate1361 ( .A(N5498), .B(N4332), .Y(N6120) );
  AND2X1 gate1362_1 ( .A(N5506), .B(N5498), .Y(N6121_1) );
  AND2X1 gate1362 ( .A(N4336), .B(N6121_1), .Y(N6121) );
  AND2X1 gate1363_1 ( .A(N5520), .B(N5498), .Y(N6122_1) );
  AND2X1 gate1363_2 ( .A(N4342), .B(N5506), .Y(N6122_2) );
  AND2X1 gate1363 ( .A(N6122_1), .B(N6122_2), .Y(N6122) );
  AND2X1 gate1364_1 ( .A(N5536), .B(N5520), .Y(N6123_1) );
  AND2X1 gate1364_2 ( .A(N5498), .B(N4349), .Y(N6123_2) );
  AND2X1 gate1364_3 ( .A(N5506), .B(N6123_1), .Y(N6123_3) );
  AND2X1 gate1364 ( .A(N6123_2), .B(N6123_3), .Y(N6123) );
  AND2X1 gate1365 ( .A(N5506), .B(N4336), .Y(N6124) );
  AND2X1 gate1366_1 ( .A(N5520), .B(N4342), .Y(N6125_1) );
  AND2X1 gate1366 ( .A(N5506), .B(N6125_1), .Y(N6125) );
  AND2X1 gate1367_1 ( .A(N5536), .B(N5520), .Y(N6126_1) );
  AND2X1 gate1367_2 ( .A(N4349), .B(N5506), .Y(N6126_2) );
  AND2X1 gate1367 ( .A(N6126_1), .B(N6126_2), .Y(N6126) );
  AND2X1 gate1368_1 ( .A(N5555), .B(N5520), .Y(N6127_1) );
  AND2X1 gate1368_2 ( .A(N5506), .B(N5536), .Y(N6127_2) );
  AND2X1 gate1368 ( .A(N6127_1), .B(N6127_2), .Y(N6127) );
  AND2X1 gate1369 ( .A(N5506), .B(N4336), .Y(N6128) );
  AND2X1 gate1370_1 ( .A(N5520), .B(N4342), .Y(N6129_1) );
  AND2X1 gate1370 ( .A(N5506), .B(N6129_1), .Y(N6129) );
  AND2X1 gate1371_1 ( .A(N5536), .B(N5520), .Y(N6130_1) );
  AND2X1 gate1371_2 ( .A(N4349), .B(N5506), .Y(N6130_2) );
  AND2X1 gate1371 ( .A(N6130_1), .B(N6130_2), .Y(N6130) );
  AND2X1 gate1372 ( .A(N5520), .B(N4342), .Y(N6131) );
  AND2X1 gate1373_1 ( .A(N5536), .B(N5520), .Y(N6132_1) );
  AND2X1 gate1373 ( .A(N4349), .B(N6132_1), .Y(N6132) );
  AND2X1 gate1374_1 ( .A(N5555), .B(N5520), .Y(N6133_1) );
  AND2X1 gate1374 ( .A(N5536), .B(N6133_1), .Y(N6133) );
  AND2X1 gate1375 ( .A(N5520), .B(N4342), .Y(N6134) );
  AND2X1 gate1376_1 ( .A(N5536), .B(N5520), .Y(N6135_1) );
  AND2X1 gate1376 ( .A(N4349), .B(N6135_1), .Y(N6135) );
  AND2X1 gate1377 ( .A(N5536), .B(N4349), .Y(N6136) );
  AND2X1 gate1378 ( .A(N5549), .B(N5488), .Y(N6137) );
  AND2X1 gate1379 ( .A(N5555), .B(N5536), .Y(N6138) );
  INVX1 gate1380 ( .A(N5573), .Y(N6139) );
  AND2X1 gate1381_1 ( .A(N4364), .B(N5573), .Y(N6140_1) );
  AND2X1 gate1381_2 ( .A(N5562), .B(N4357), .Y(N6140_2) );
  AND2X1 gate1381 ( .A(N6140_1), .B(N6140_2), .Y(N6140) );
  AND2X1 gate1382_1 ( .A(N5562), .B(N4385), .Y(N6143_1) );
  AND2X1 gate1382 ( .A(N4364), .B(N6143_1), .Y(N6143) );
  AND2X1 gate1383_1 ( .A(N5573), .B(N5562), .Y(N6144_1) );
  AND2X1 gate1383 ( .A(N4364), .B(N6144_1), .Y(N6144) );
  AND2X1 gate1384_1 ( .A(N4385), .B(N5562), .Y(N6145_1) );
  AND2X1 gate1384 ( .A(N4364), .B(N6145_1), .Y(N6145) );
  AND2X1 gate1385 ( .A(N5562), .B(N4385), .Y(N6146) );
  AND2X1 gate1386 ( .A(N5573), .B(N5562), .Y(N6147) );
  AND2X1 gate1387 ( .A(N5562), .B(N4385), .Y(N6148) );
  AND2X1 gate1388_1 ( .A(N5264), .B(N4405), .Y(N6149_1) );
  AND2X1 gate1388_2 ( .A(N5595), .B(N5579), .Y(N6149_2) );
  AND2X1 gate1388_3 ( .A(N5606), .B(N6149_1), .Y(N6149_3) );
  AND2X1 gate1388 ( .A(N6149_2), .B(N6149_3), .Y(N6149) );
  AND2X1 gate1389 ( .A(N5579), .B(N4067), .Y(N6152) );
  AND2X1 gate1390_1 ( .A(N5264), .B(N5579), .Y(N6153_1) );
  AND2X1 gate1390 ( .A(N4396), .B(N6153_1), .Y(N6153) );
  AND2X1 gate1391_1 ( .A(N5595), .B(N5579), .Y(N6154_1) );
  AND2X1 gate1391_2 ( .A(N4400), .B(N5264), .Y(N6154_2) );
  AND2X1 gate1391 ( .A(N6154_1), .B(N6154_2), .Y(N6154) );
  AND2X1 gate1392_1 ( .A(N5606), .B(N5595), .Y(N6155_1) );
  AND2X1 gate1392_2 ( .A(N5579), .B(N4412), .Y(N6155_2) );
  AND2X1 gate1392_3 ( .A(N5264), .B(N6155_1), .Y(N6155_3) );
  AND2X1 gate1392 ( .A(N6155_2), .B(N6155_3), .Y(N6155) );
  AND2X1 gate1393_1 ( .A(N5595), .B(N4400), .Y(N6156_1) );
  AND2X1 gate1393 ( .A(N5264), .B(N6156_1), .Y(N6156) );
  AND2X1 gate1394_1 ( .A(N5606), .B(N5595), .Y(N6157_1) );
  AND2X1 gate1394_2 ( .A(N4412), .B(N5264), .Y(N6157_2) );
  AND2X1 gate1394 ( .A(N6157_1), .B(N6157_2), .Y(N6157) );
  AND2X1 gate1395_1 ( .A(N54), .B(N4405), .Y(N6158_1) );
  AND2X1 gate1395_2 ( .A(N5595), .B(N5606), .Y(N6158_2) );
  AND2X1 gate1395_3 ( .A(N5264), .B(N6158_1), .Y(N6158_3) );
  AND2X1 gate1395 ( .A(N6158_2), .B(N6158_3), .Y(N6158) );
  AND2X1 gate1396 ( .A(N4400), .B(N5595), .Y(N6159) );
  AND2X1 gate1397_1 ( .A(N5606), .B(N5595), .Y(N6160_1) );
  AND2X1 gate1397 ( .A(N4412), .B(N6160_1), .Y(N6160) );
  AND2X1 gate1398_1 ( .A(N54), .B(N4405), .Y(N6161_1) );
  AND2X1 gate1398_2 ( .A(N5595), .B(N5606), .Y(N6161_2) );
  AND2X1 gate1398 ( .A(N6161_1), .B(N6161_2), .Y(N6161) );
  AND2X1 gate1399 ( .A(N5606), .B(N4412), .Y(N6162) );
  AND2X1 gate1400_1 ( .A(N54), .B(N4405), .Y(N6163_1) );
  AND2X1 gate1400 ( .A(N5606), .B(N6163_1), .Y(N6163) );
  NAND2X1 gate1401 ( .A(N5616), .B(N5955), .Y(N6164) );
  AND2X1 gate1402_1 ( .A(N5684), .B(N5624), .Y(N6168_1) );
  AND2X1 gate1402_2 ( .A(N4425), .B(N4418), .Y(N6168_2) );
  AND2X1 gate1402 ( .A(N6168_1), .B(N6168_2), .Y(N6168) );
  AND2X1 gate1403_1 ( .A(N5624), .B(N4445), .Y(N6171_1) );
  AND2X1 gate1403 ( .A(N4425), .B(N6171_1), .Y(N6171) );
  AND2X1 gate1404_1 ( .A(N5684), .B(N5624), .Y(N6172_1) );
  AND2X1 gate1404 ( .A(N4425), .B(N6172_1), .Y(N6172) );
  AND2X1 gate1405_1 ( .A(N5624), .B(N4445), .Y(N6173_1) );
  AND2X1 gate1405 ( .A(N4425), .B(N6173_1), .Y(N6173) );
  AND2X1 gate1406 ( .A(N5624), .B(N4445), .Y(N6174) );
  AND2X1 gate1407_1 ( .A(N4477), .B(N5671), .Y(N6175_1) );
  AND2X1 gate1407_2 ( .A(N5655), .B(N5284), .Y(N6175_2) );
  AND2X1 gate1407_3 ( .A(N5634), .B(N6175_1), .Y(N6175_3) );
  AND2X1 gate1407 ( .A(N6175_2), .B(N6175_3), .Y(N6175) );
  AND2X1 gate1408 ( .A(N5634), .B(N4080), .Y(N6178) );
  AND2X1 gate1409_1 ( .A(N5284), .B(N5634), .Y(N6179_1) );
  AND2X1 gate1409 ( .A(N4456), .B(N6179_1), .Y(N6179) );
  AND2X1 gate1410_1 ( .A(N5655), .B(N5634), .Y(N6180_1) );
  AND2X1 gate1410_2 ( .A(N4462), .B(N5284), .Y(N6180_2) );
  AND2X1 gate1410 ( .A(N6180_1), .B(N6180_2), .Y(N6180) );
  AND2X1 gate1411_1 ( .A(N5671), .B(N5655), .Y(N6181_1) );
  AND2X1 gate1411_2 ( .A(N5634), .B(N4469), .Y(N6181_2) );
  AND2X1 gate1411_3 ( .A(N5284), .B(N6181_1), .Y(N6181_3) );
  AND2X1 gate1411 ( .A(N6181_2), .B(N6181_3), .Y(N6181) );
  AND2X1 gate1412_1 ( .A(N5655), .B(N4462), .Y(N6182_1) );
  AND2X1 gate1412 ( .A(N5284), .B(N6182_1), .Y(N6182) );
  AND2X1 gate1413_1 ( .A(N5671), .B(N5655), .Y(N6183_1) );
  AND2X1 gate1413_2 ( .A(N4469), .B(N5284), .Y(N6183_2) );
  AND2X1 gate1413 ( .A(N6183_1), .B(N6183_2), .Y(N6183) );
  AND2X1 gate1414_1 ( .A(N4477), .B(N5655), .Y(N6184_1) );
  AND2X1 gate1414_2 ( .A(N5284), .B(N5671), .Y(N6184_2) );
  AND2X1 gate1414 ( .A(N6184_1), .B(N6184_2), .Y(N6184) );
  AND2X1 gate1415_1 ( .A(N5655), .B(N4462), .Y(N6185_1) );
  AND2X1 gate1415 ( .A(N5284), .B(N6185_1), .Y(N6185) );
  AND2X1 gate1416_1 ( .A(N5671), .B(N5655), .Y(N6186_1) );
  AND2X1 gate1416_2 ( .A(N4469), .B(N5284), .Y(N6186_2) );
  AND2X1 gate1416 ( .A(N6186_1), .B(N6186_2), .Y(N6186) );
  AND2X1 gate1417 ( .A(N5655), .B(N4462), .Y(N6187) );
  AND2X1 gate1418_1 ( .A(N5671), .B(N5655), .Y(N6188_1) );
  AND2X1 gate1418 ( .A(N4469), .B(N6188_1), .Y(N6188) );
  AND2X1 gate1419_1 ( .A(N4477), .B(N5655), .Y(N6189_1) );
  AND2X1 gate1419 ( .A(N5671), .B(N6189_1), .Y(N6189) );
  AND2X1 gate1420 ( .A(N5655), .B(N4462), .Y(N6190) );
  AND2X1 gate1421_1 ( .A(N5671), .B(N5655), .Y(N6191_1) );
  AND2X1 gate1421 ( .A(N4469), .B(N6191_1), .Y(N6191) );
  AND2X1 gate1422 ( .A(N5671), .B(N4469), .Y(N6192) );
  AND2X1 gate1423 ( .A(N5684), .B(N5624), .Y(N6193) );
  AND2X1 gate1424 ( .A(N4477), .B(N5671), .Y(N6194) );
  INVX1 gate1425 ( .A(N5692), .Y(N6197) );
  INVX1 gate1426 ( .A(N5696), .Y(N6200) );
  INVX1 gate1427 ( .A(N5703), .Y(N6203) );
  INVX1 gate1428 ( .A(N5707), .Y(N6206) );
  BUFX2 gate1429 ( .A(N5700), .Y(N6209) );
  BUFX2 gate1430 ( .A(N5700), .Y(N6212) );
  BUFX2 gate1431 ( .A(N5711), .Y(N6215) );
  BUFX2 gate1432 ( .A(N5711), .Y(N6218) );
  NAND2X1 gate1433 ( .A(N5049), .B(N6023), .Y(N6221) );
  INVX1 gate1434 ( .A(N5756), .Y(N6234) );
  NAND2X1 gate1435 ( .A(N5756), .B(N6044), .Y(N6235) );
  BUFX2 gate1436 ( .A(N5462), .Y(N6238) );
  BUFX2 gate1437 ( .A(N5389), .Y(N6241) );
  BUFX2 gate1438 ( .A(N5389), .Y(N6244) );
  BUFX2 gate1439 ( .A(N5396), .Y(N6247) );
  BUFX2 gate1440 ( .A(N5396), .Y(N6250) );
  BUFX2 gate1441 ( .A(N5407), .Y(N6253) );
  BUFX2 gate1442 ( .A(N5407), .Y(N6256) );
  BUFX2 gate1443 ( .A(N5424), .Y(N6259) );
  BUFX2 gate1444 ( .A(N5431), .Y(N6262) );
  BUFX2 gate1445 ( .A(N5441), .Y(N6265) );
  BUFX2 gate1446 ( .A(N5452), .Y(N6268) );
  BUFX2 gate1447 ( .A(N5549), .Y(N6271) );
  BUFX2 gate1448 ( .A(N5488), .Y(N6274) );
  BUFX2 gate1449 ( .A(N5470), .Y(N6277) );
  BUFX2 gate1450 ( .A(N5477), .Y(N6280) );
  BUFX2 gate1451 ( .A(N5549), .Y(N6283) );
  BUFX2 gate1452 ( .A(N5488), .Y(N6286) );
  BUFX2 gate1453 ( .A(N5470), .Y(N6289) );
  BUFX2 gate1454 ( .A(N5477), .Y(N6292) );
  BUFX2 gate1455 ( .A(N5555), .Y(N6295) );
  BUFX2 gate1456 ( .A(N5536), .Y(N6298) );
  BUFX2 gate1457 ( .A(N5498), .Y(N6301) );
  BUFX2 gate1458 ( .A(N5520), .Y(N6304) );
  BUFX2 gate1459 ( .A(N5506), .Y(N6307) );
  BUFX2 gate1460 ( .A(N5506), .Y(N6310) );
  BUFX2 gate1461 ( .A(N5555), .Y(N6313) );
  BUFX2 gate1462 ( .A(N5536), .Y(N6316) );
  BUFX2 gate1463 ( .A(N5498), .Y(N6319) );
  BUFX2 gate1464 ( .A(N5520), .Y(N6322) );
  BUFX2 gate1465 ( .A(N5562), .Y(N6325) );
  BUFX2 gate1466 ( .A(N5562), .Y(N6328) );
  BUFX2 gate1467 ( .A(N5579), .Y(N6331) );
  BUFX2 gate1468 ( .A(N5595), .Y(N6335) );
  BUFX2 gate1469 ( .A(N5606), .Y(N6338) );
  BUFX2 gate1470 ( .A(N5684), .Y(N6341) );
  BUFX2 gate1471 ( .A(N5624), .Y(N6344) );
  BUFX2 gate1472 ( .A(N5684), .Y(N6347) );
  BUFX2 gate1473 ( .A(N5624), .Y(N6350) );
  BUFX2 gate1474 ( .A(N5671), .Y(N6353) );
  BUFX2 gate1475 ( .A(N5634), .Y(N6356) );
  BUFX2 gate1476 ( .A(N5655), .Y(N6359) );
  BUFX2 gate1477 ( .A(N5671), .Y(N6364) );
  BUFX2 gate1478 ( .A(N5634), .Y(N6367) );
  BUFX2 gate1479 ( .A(N5655), .Y(N6370) );
  INVX1 gate1480 ( .A(N5736), .Y(N6373) );
  INVX1 gate1481 ( .A(N5739), .Y(N6374) );
  INVX1 gate1482 ( .A(N5742), .Y(N6375) );
  INVX1 gate1483 ( .A(N5745), .Y(N6376) );
  NAND2X1 gate1484 ( .A(N4243), .B(N6065), .Y(N6377) );
  NAND2X1 gate1485 ( .A(N5236), .B(N6068), .Y(N6378) );
  OR2X1 gate1486_1 ( .A(N4268), .B(N6071), .Y(N6382_1) );
  OR2X1 gate1486_2 ( .A(N6072), .B(N6073), .Y(N6382_2) );
  OR2X1 gate1486 ( .A(N6382_1), .B(N6382_2), .Y(N6382) );
  OR2X1 gate1487_1 ( .A(N3968), .B(N5065), .Y(N6386_1) );
  OR2X1 gate1487_2 ( .A(N5066), .B(N6074), .Y(N6386_2) );
  OR2X1 gate1487 ( .A(N6386_1), .B(N6386_2), .Y(N6386) );
  OR2X1 gate1488_1 ( .A(N4271), .B(N6075), .Y(N6388_1) );
  OR2X1 gate1488_2 ( .A(N6076), .B(N6077), .Y(N6388_2) );
  OR2X1 gate1488 ( .A(N6388_1), .B(N6388_2), .Y(N6388) );
  OR2X1 gate1489_1 ( .A(N3968), .B(N5067), .Y(N6392_1) );
  OR2X1 gate1489_2 ( .A(N5068), .B(N6078), .Y(N6392_2) );
  OR2X1 gate1489 ( .A(N6392_1), .B(N6392_2), .Y(N6392) );
  OR2X1 gate1490_1 ( .A(N4297), .B(N6094), .Y(N6397_1) );
  OR2X1 gate1490_2 ( .A(N6095), .B(N6096), .Y(N6397_2) );
  OR2X1 gate1490_3 ( .A(N6097), .B(N6397_1), .Y(N6397_3) );
  OR2X1 gate1490 ( .A(N6397_2), .B(N6397_3), .Y(N6397) );
  OR2X1 gate1491 ( .A(N4320), .B(N6116), .Y(N6411) );
  OR2X1 gate1492_1 ( .A(N4331), .B(N6120), .Y(N6415_1) );
  OR2X1 gate1492_2 ( .A(N6121), .B(N6122), .Y(N6415_2) );
  OR2X1 gate1492_3 ( .A(N6123), .B(N6415_1), .Y(N6415_3) );
  OR2X1 gate1492 ( .A(N6415_2), .B(N6415_3), .Y(N6415) );
  OR2X1 gate1493 ( .A(N4342), .B(N6136), .Y(N6419) );
  OR2X1 gate1494_1 ( .A(N4392), .B(N6152), .Y(N6427_1) );
  OR2X1 gate1494_2 ( .A(N6153), .B(N6154), .Y(N6427_2) );
  OR2X1 gate1494_3 ( .A(N6155), .B(N6427_1), .Y(N6427_3) );
  OR2X1 gate1494 ( .A(N6427_2), .B(N6427_3), .Y(N6427) );
  INVX1 gate1495 ( .A(N6048), .Y(N6434) );
  OR2X1 gate1496 ( .A(N4440), .B(N6174), .Y(N6437) );
  OR2X1 gate1497_1 ( .A(N4451), .B(N6178), .Y(N6441_1) );
  OR2X1 gate1497_2 ( .A(N6179), .B(N6180), .Y(N6441_2) );
  OR2X1 gate1497_3 ( .A(N6181), .B(N6441_1), .Y(N6441_3) );
  OR2X1 gate1497 ( .A(N6441_2), .B(N6441_3), .Y(N6441) );
  OR2X1 gate1498 ( .A(N4462), .B(N6192), .Y(N6445) );
  INVX1 gate1499 ( .A(N6051), .Y(N6448) );
  INVX1 gate1500 ( .A(N6054), .Y(N6449) );
  NAND2X1 gate1501 ( .A(N6221), .B(N6024), .Y(N6466) );
  INVX1 gate1502 ( .A(N6031), .Y(N6469) );
  INVX1 gate1503 ( .A(N6034), .Y(N6470) );
  INVX1 gate1504 ( .A(N6037), .Y(N6471) );
  INVX1 gate1505 ( .A(N6040), .Y(N6472) );
  AND2X1 gate1506_1 ( .A(N5315), .B(N4524), .Y(N6473_1) );
  AND2X1 gate1506 ( .A(N6031), .B(N6473_1), .Y(N6473) );
  AND2X1 gate1507_1 ( .A(N6025), .B(N5150), .Y(N6474_1) );
  AND2X1 gate1507 ( .A(N6034), .B(N6474_1), .Y(N6474) );
  AND2X1 gate1508_1 ( .A(N5324), .B(N4532), .Y(N6475_1) );
  AND2X1 gate1508 ( .A(N6037), .B(N6475_1), .Y(N6475) );
  AND2X1 gate1509_1 ( .A(N6028), .B(N5157), .Y(N6476_1) );
  AND2X1 gate1509 ( .A(N6040), .B(N6476_1), .Y(N6476) );
  NAND2X1 gate1510 ( .A(N5385), .B(N6234), .Y(N6477) );
  NAND2X1 gate1511 ( .A(N6045), .B(N132), .Y(N6478) );
  OR2X1 gate1512_1 ( .A(N4280), .B(N6083), .Y(N6482_1) );
  OR2X1 gate1512_2 ( .A(N6084), .B(N6085), .Y(N6482_2) );
  OR2X1 gate1512 ( .A(N6482_1), .B(N6482_2), .Y(N6482) );
  NOR3X1 gate1513 ( .A(N4280), .B(N6086), .C(N6087), .Y(N6486) );
  OR2X1 gate1514_1 ( .A(N4284), .B(N6088), .Y(N6490_1) );
  OR2X1 gate1514 ( .A(N6089), .B(N6490_1), .Y(N6490) );
  NOR2X1 gate1515 ( .A(N4284), .B(N6090), .Y(N6494) );
  OR2X1 gate1516_1 ( .A(N4298), .B(N6098), .Y(N6500_1) );
  OR2X1 gate1516_2 ( .A(N6099), .B(N6100), .Y(N6500_2) );
  OR2X1 gate1516_3 ( .A(N6101), .B(N6500_1), .Y(N6500_3) );
  OR2X1 gate1516 ( .A(N6500_2), .B(N6500_3), .Y(N6500) );
  OR2X1 gate1517_1 ( .A(N4301), .B(N6102), .Y(N6504_1) );
  OR2X1 gate1517_2 ( .A(N6103), .B(N6104), .Y(N6504_2) );
  OR2X1 gate1517 ( .A(N6504_1), .B(N6504_2), .Y(N6504) );
  OR2X1 gate1518_1 ( .A(N4305), .B(N6105), .Y(N6508_1) );
  OR2X1 gate1518 ( .A(N6106), .B(N6508_1), .Y(N6508) );
  OR2X1 gate1519 ( .A(N4310), .B(N6107), .Y(N6512) );
  OR2X1 gate1520_1 ( .A(N4316), .B(N6111), .Y(N6516_1) );
  OR2X1 gate1520_2 ( .A(N6112), .B(N6113), .Y(N6516_2) );
  OR2X1 gate1520 ( .A(N6516_1), .B(N6516_2), .Y(N6516) );
  NOR3X1 gate1521 ( .A(N4316), .B(N6114), .C(N6115), .Y(N6526) );
  OR2X1 gate1522_1 ( .A(N4336), .B(N6131), .Y(N6536_1) );
  OR2X1 gate1522_2 ( .A(N6132), .B(N6133), .Y(N6536_2) );
  OR2X1 gate1522 ( .A(N6536_1), .B(N6536_2), .Y(N6536) );
  OR2X1 gate1523_1 ( .A(N4332), .B(N6124), .Y(N6539_1) );
  OR2X1 gate1523_2 ( .A(N6125), .B(N6126), .Y(N6539_2) );
  OR2X1 gate1523_3 ( .A(N6127), .B(N6539_1), .Y(N6539_3) );
  OR2X1 gate1523 ( .A(N6539_2), .B(N6539_3), .Y(N6539) );
  NOR3X1 gate1524 ( .A(N4336), .B(N6134), .C(N6135), .Y(N6553) );
  NOR2X1 gate1525_1 ( .A(N4332), .B(N6128), .Y(N6556_1) );
  NOR2X1 gate1525_2 ( .A(N6129), .B(N6130), .Y(N6556_2) );
  NOR2X1 gate1525 ( .A(N6556_1), .B(N6556_2), .Y(N6556) );
  OR2X1 gate1526_1 ( .A(N4375), .B(N5117), .Y(N6566_1) );
  OR2X1 gate1526_2 ( .A(N6143), .B(N6144), .Y(N6566_2) );
  OR2X1 gate1526 ( .A(N6566_1), .B(N6566_2), .Y(N6566) );
  NOR3X1 gate1527 ( .A(N4375), .B(N5118), .C(N6145), .Y(N6569) );
  OR2X1 gate1528_1 ( .A(N4379), .B(N6146), .Y(N6572_1) );
  OR2X1 gate1528 ( .A(N6147), .B(N6572_1), .Y(N6572) );
  NOR2X1 gate1529 ( .A(N4379), .B(N6148), .Y(N6575) );
  OR2X1 gate1530_1 ( .A(N4067), .B(N5954), .Y(N6580_1) );
  OR2X1 gate1530_2 ( .A(N6156), .B(N6157), .Y(N6580_2) );
  OR2X1 gate1530_3 ( .A(N6158), .B(N6580_1), .Y(N6580_3) );
  OR2X1 gate1530 ( .A(N6580_2), .B(N6580_3), .Y(N6580) );
  OR2X1 gate1531_1 ( .A(N4396), .B(N6159), .Y(N6584_1) );
  OR2X1 gate1531_2 ( .A(N6160), .B(N6161), .Y(N6584_2) );
  OR2X1 gate1531 ( .A(N6584_1), .B(N6584_2), .Y(N6584) );
  OR2X1 gate1532_1 ( .A(N4400), .B(N6162), .Y(N6587_1) );
  OR2X1 gate1532 ( .A(N6163), .B(N6587_1), .Y(N6587) );
  OR2X1 gate1533_1 ( .A(N4436), .B(N5132), .Y(N6592_1) );
  OR2X1 gate1533_2 ( .A(N6171), .B(N6172), .Y(N6592_2) );
  OR2X1 gate1533 ( .A(N6592_1), .B(N6592_2), .Y(N6592) );
  NOR3X1 gate1534 ( .A(N4436), .B(N5133), .C(N6173), .Y(N6599) );
  OR2X1 gate1535_1 ( .A(N4456), .B(N6187), .Y(N6606_1) );
  OR2X1 gate1535_2 ( .A(N6188), .B(N6189), .Y(N6606_2) );
  OR2X1 gate1535 ( .A(N6606_1), .B(N6606_2), .Y(N6606) );
  OR2X1 gate1536_1 ( .A(N4080), .B(N6005), .Y(N6609_1) );
  OR2X1 gate1536_2 ( .A(N6182), .B(N6183), .Y(N6609_2) );
  OR2X1 gate1536_3 ( .A(N6184), .B(N6609_1), .Y(N6609_3) );
  OR2X1 gate1536 ( .A(N6609_2), .B(N6609_3), .Y(N6609) );
  NOR3X1 gate1537 ( .A(N4456), .B(N6190), .C(N6191), .Y(N6619) );
  NOR2X1 gate1538_1 ( .A(N4080), .B(N6006), .Y(N6622_1) );
  NOR2X1 gate1538_2 ( .A(N6185), .B(N6186), .Y(N6622_2) );
  NOR2X1 gate1538 ( .A(N6622_1), .B(N6622_2), .Y(N6622) );
  NAND2X1 gate1539 ( .A(N5739), .B(N6373), .Y(N6630) );
  NAND2X1 gate1540 ( .A(N5736), .B(N6374), .Y(N6631) );
  NAND2X1 gate1541 ( .A(N5745), .B(N6375), .Y(N6632) );
  NAND2X1 gate1542 ( .A(N5742), .B(N6376), .Y(N6633) );
  NAND2X1 gate1543 ( .A(N6377), .B(N6066), .Y(N6634) );
  NAND2X1 gate1544 ( .A(N6069), .B(N6378), .Y(N6637) );
  INVX1 gate1545 ( .A(N6164), .Y(N6640) );
  AND2X1 gate1546 ( .A(N6108), .B(N6117), .Y(N6641) );
  AND2X1 gate1547 ( .A(N6140), .B(N6149), .Y(N6643) );
  AND2X1 gate1548 ( .A(N6168), .B(N6175), .Y(N6646) );
  AND2X1 gate1549 ( .A(N6080), .B(N6091), .Y(N6648) );
  NAND2X1 gate1550 ( .A(N6238), .B(N2637), .Y(N6650) );
  INVX1 gate1551 ( .A(N6238), .Y(N6651) );
  INVX1 gate1552 ( .A(N6241), .Y(N6653) );
  INVX1 gate1553 ( .A(N6244), .Y(N6655) );
  INVX1 gate1554 ( .A(N6247), .Y(N6657) );
  INVX1 gate1555 ( .A(N6250), .Y(N6659) );
  NAND2X1 gate1556 ( .A(N6253), .B(N5087), .Y(N6660) );
  INVX1 gate1557 ( .A(N6253), .Y(N6661) );
  NAND2X1 gate1558 ( .A(N6256), .B(N5469), .Y(N6662) );
  INVX1 gate1559 ( .A(N6256), .Y(N6663) );
  AND2X1 gate1560 ( .A(N6091), .B(N4), .Y(N6664) );
  INVX1 gate1561 ( .A(N6259), .Y(N6666) );
  INVX1 gate1562 ( .A(N6262), .Y(N6668) );
  INVX1 gate1563 ( .A(N6265), .Y(N6670) );
  INVX1 gate1564 ( .A(N6268), .Y(N6672) );
  INVX1 gate1565 ( .A(N6117), .Y(N6675) );
  INVX1 gate1566 ( .A(N6280), .Y(N6680) );
  INVX1 gate1567 ( .A(N6292), .Y(N6681) );
  INVX1 gate1568 ( .A(N6307), .Y(N6682) );
  INVX1 gate1569 ( .A(N6310), .Y(N6683) );
  NAND2X1 gate1570 ( .A(N6325), .B(N5120), .Y(N6689) );
  INVX1 gate1571 ( .A(N6325), .Y(N6690) );
  NAND2X1 gate1572 ( .A(N6328), .B(N5622), .Y(N6691) );
  INVX1 gate1573 ( .A(N6328), .Y(N6692) );
  AND2X1 gate1574 ( .A(N6149), .B(N54), .Y(N6693) );
  INVX1 gate1575 ( .A(N6331), .Y(N6695) );
  INVX1 gate1576 ( .A(N6335), .Y(N6698) );
  NAND2X1 gate1577 ( .A(N6338), .B(N5956), .Y(N6699) );
  INVX1 gate1578 ( .A(N6338), .Y(N6700) );
  INVX1 gate1579 ( .A(N6175), .Y(N6703) );
  INVX1 gate1580 ( .A(N6209), .Y(N6708) );
  INVX1 gate1581 ( .A(N6212), .Y(N6709) );
  INVX1 gate1582 ( .A(N6215), .Y(N6710) );
  INVX1 gate1583 ( .A(N6218), .Y(N6711) );
  AND2X1 gate1584_1 ( .A(N5696), .B(N5692), .Y(N6712_1) );
  AND2X1 gate1584 ( .A(N6209), .B(N6712_1), .Y(N6712) );
  AND2X1 gate1585_1 ( .A(N6200), .B(N6197), .Y(N6713_1) );
  AND2X1 gate1585 ( .A(N6212), .B(N6713_1), .Y(N6713) );
  AND2X1 gate1586_1 ( .A(N5707), .B(N5703), .Y(N6714_1) );
  AND2X1 gate1586 ( .A(N6215), .B(N6714_1), .Y(N6714) );
  AND2X1 gate1587_1 ( .A(N6206), .B(N6203), .Y(N6715_1) );
  AND2X1 gate1587 ( .A(N6218), .B(N6715_1), .Y(N6715) );
  BUFX2 gate1588 ( .A(N6466), .Y(N6716) );
  AND2X1 gate1589_1 ( .A(N6164), .B(N1777), .Y(N6718_1) );
  AND2X1 gate1589 ( .A(N3130), .B(N6718_1), .Y(N6718) );
  AND2X1 gate1590_1 ( .A(N5150), .B(N5315), .Y(N6719_1) );
  AND2X1 gate1590 ( .A(N6469), .B(N6719_1), .Y(N6719) );
  AND2X1 gate1591_1 ( .A(N4524), .B(N6025), .Y(N6720_1) );
  AND2X1 gate1591 ( .A(N6470), .B(N6720_1), .Y(N6720) );
  AND2X1 gate1592_1 ( .A(N5157), .B(N5324), .Y(N6721_1) );
  AND2X1 gate1592 ( .A(N6471), .B(N6721_1), .Y(N6721) );
  AND2X1 gate1593_1 ( .A(N4532), .B(N6028), .Y(N6722_1) );
  AND2X1 gate1593 ( .A(N6472), .B(N6722_1), .Y(N6722) );
  NAND2X1 gate1594 ( .A(N6477), .B(N6235), .Y(N6724) );
  INVX1 gate1595 ( .A(N6271), .Y(N6739) );
  INVX1 gate1596 ( .A(N6274), .Y(N6740) );
  INVX1 gate1597 ( .A(N6277), .Y(N6741) );
  INVX1 gate1598 ( .A(N6283), .Y(N6744) );
  INVX1 gate1599 ( .A(N6286), .Y(N6745) );
  INVX1 gate1600 ( .A(N6289), .Y(N6746) );
  INVX1 gate1601 ( .A(N6295), .Y(N6751) );
  INVX1 gate1602 ( .A(N6298), .Y(N6752) );
  INVX1 gate1603 ( .A(N6301), .Y(N6753) );
  INVX1 gate1604 ( .A(N6304), .Y(N6754) );
  INVX1 gate1605 ( .A(N6322), .Y(N6755) );
  INVX1 gate1606 ( .A(N6313), .Y(N6760) );
  INVX1 gate1607 ( .A(N6316), .Y(N6761) );
  INVX1 gate1608 ( .A(N6319), .Y(N6762) );
  INVX1 gate1609 ( .A(N6341), .Y(N6772) );
  INVX1 gate1610 ( .A(N6344), .Y(N6773) );
  INVX1 gate1611 ( .A(N6347), .Y(N6776) );
  INVX1 gate1612 ( .A(N6350), .Y(N6777) );
  INVX1 gate1613 ( .A(N6353), .Y(N6782) );
  INVX1 gate1614 ( .A(N6356), .Y(N6783) );
  INVX1 gate1615 ( .A(N6359), .Y(N6784) );
  INVX1 gate1616 ( .A(N6370), .Y(N6785) );
  INVX1 gate1617 ( .A(N6364), .Y(N6790) );
  INVX1 gate1618 ( .A(N6367), .Y(N6791) );
  NAND2X1 gate1619 ( .A(N6630), .B(N6631), .Y(N6792) );
  NAND2X1 gate1620 ( .A(N6632), .B(N6633), .Y(N6795) );
  AND2X1 gate1621 ( .A(N6108), .B(N6415), .Y(N6801) );
  AND2X1 gate1622 ( .A(N6427), .B(N6140), .Y(N6802) );
  AND2X1 gate1623 ( .A(N6397), .B(N6080), .Y(N6803) );
  AND2X1 gate1624 ( .A(N6168), .B(N6441), .Y(N6804) );
  INVX1 gate1625 ( .A(N6466), .Y(N6805) );
  NAND2X1 gate1626 ( .A(N1851), .B(N6651), .Y(N6806) );
  INVX1 gate1627 ( .A(N6482), .Y(N6807) );
  NAND2X1 gate1628 ( .A(N6482), .B(N6653), .Y(N6808) );
  INVX1 gate1629 ( .A(N6486), .Y(N6809) );
  NAND2X1 gate1630 ( .A(N6486), .B(N6655), .Y(N6810) );
  INVX1 gate1631 ( .A(N6490), .Y(N6811) );
  NAND2X1 gate1632 ( .A(N6490), .B(N6657), .Y(N6812) );
  INVX1 gate1633 ( .A(N6494), .Y(N6813) );
  NAND2X1 gate1634 ( .A(N6494), .B(N6659), .Y(N6814) );
  NAND2X1 gate1635 ( .A(N4575), .B(N6661), .Y(N6815) );
  NAND2X1 gate1636 ( .A(N5169), .B(N6663), .Y(N6816) );
  OR2X1 gate1637 ( .A(N6397), .B(N6664), .Y(N6817) );
  INVX1 gate1638 ( .A(N6500), .Y(N6823) );
  NAND2X1 gate1639 ( .A(N6500), .B(N6666), .Y(N6824) );
  INVX1 gate1640 ( .A(N6504), .Y(N6825) );
  NAND2X1 gate1641 ( .A(N6504), .B(N6668), .Y(N6826) );
  INVX1 gate1642 ( .A(N6508), .Y(N6827) );
  NAND2X1 gate1643 ( .A(N6508), .B(N6670), .Y(N6828) );
  INVX1 gate1644 ( .A(N6512), .Y(N6829) );
  NAND2X1 gate1645 ( .A(N6512), .B(N6672), .Y(N6830) );
  INVX1 gate1646 ( .A(N6415), .Y(N6831) );
  INVX1 gate1647 ( .A(N6566), .Y(N6834) );
  NAND2X1 gate1648 ( .A(N6566), .B(N5618), .Y(N6835) );
  INVX1 gate1649 ( .A(N6569), .Y(N6836) );
  NAND2X1 gate1650 ( .A(N6569), .B(N5619), .Y(N6837) );
  INVX1 gate1651 ( .A(N6572), .Y(N6838) );
  NAND2X1 gate1652 ( .A(N6572), .B(N5620), .Y(N6839) );
  INVX1 gate1653 ( .A(N6575), .Y(N6840) );
  NAND2X1 gate1654 ( .A(N6575), .B(N5621), .Y(N6841) );
  NAND2X1 gate1655 ( .A(N4627), .B(N6690), .Y(N6842) );
  NAND2X1 gate1656 ( .A(N5195), .B(N6692), .Y(N6843) );
  OR2X1 gate1657 ( .A(N6427), .B(N6693), .Y(N6844) );
  INVX1 gate1658 ( .A(N6580), .Y(N6850) );
  NAND2X1 gate1659 ( .A(N6580), .B(N6695), .Y(N6851) );
  INVX1 gate1660 ( .A(N6584), .Y(N6852) );
  NAND2X1 gate1661 ( .A(N6584), .B(N6434), .Y(N6853) );
  INVX1 gate1662 ( .A(N6587), .Y(N6854) );
  NAND2X1 gate1663 ( .A(N6587), .B(N6698), .Y(N6855) );
  NAND2X1 gate1664 ( .A(N5346), .B(N6700), .Y(N6856) );
  INVX1 gate1665 ( .A(N6441), .Y(N6857) );
  AND2X1 gate1666_1 ( .A(N6197), .B(N5696), .Y(N6860_1) );
  AND2X1 gate1666 ( .A(N6708), .B(N6860_1), .Y(N6860) );
  AND2X1 gate1667_1 ( .A(N5692), .B(N6200), .Y(N6861_1) );
  AND2X1 gate1667 ( .A(N6709), .B(N6861_1), .Y(N6861) );
  AND2X1 gate1668_1 ( .A(N6203), .B(N5707), .Y(N6862_1) );
  AND2X1 gate1668 ( .A(N6710), .B(N6862_1), .Y(N6862) );
  AND2X1 gate1669_1 ( .A(N5703), .B(N6206), .Y(N6863_1) );
  AND2X1 gate1669 ( .A(N6711), .B(N6863_1), .Y(N6863) );
  OR2X1 gate1670_1 ( .A(N4197), .B(N6718), .Y(N6866_1) );
  OR2X1 gate1670 ( .A(N3785), .B(N6866_1), .Y(N6866) );
  NOR2X1 gate1671 ( .A(N6719), .B(N6473), .Y(N6872) );
  NOR2X1 gate1672 ( .A(N6720), .B(N6474), .Y(N6873) );
  NOR2X1 gate1673 ( .A(N6721), .B(N6475), .Y(N6874) );
  NOR2X1 gate1674 ( .A(N6722), .B(N6476), .Y(N6875) );
  INVX1 gate1675 ( .A(N6637), .Y(N6876) );
  BUFX2 gate1676 ( .A(N6724), .Y(N6877) );
  AND2X1 gate1677 ( .A(N6045), .B(N6478), .Y(N6879) );
  AND2X1 gate1678 ( .A(N6478), .B(N132), .Y(N6880) );
  OR2X1 gate1679 ( .A(N6411), .B(N6137), .Y(N6881) );
  INVX1 gate1680 ( .A(N6516), .Y(N6884) );
  INVX1 gate1681 ( .A(N6411), .Y(N6885) );
  INVX1 gate1682 ( .A(N6526), .Y(N6888) );
  INVX1 gate1683 ( .A(N6536), .Y(N6889) );
  NAND2X1 gate1684 ( .A(N6536), .B(N5176), .Y(N6890) );
  OR2X1 gate1685 ( .A(N6419), .B(N6138), .Y(N6891) );
  INVX1 gate1686 ( .A(N6539), .Y(N6894) );
  INVX1 gate1687 ( .A(N6553), .Y(N6895) );
  NAND2X1 gate1688 ( .A(N6553), .B(N5728), .Y(N6896) );
  INVX1 gate1689 ( .A(N6419), .Y(N6897) );
  INVX1 gate1690 ( .A(N6556), .Y(N6900) );
  OR2X1 gate1691 ( .A(N6437), .B(N6193), .Y(N6901) );
  INVX1 gate1692 ( .A(N6592), .Y(N6904) );
  INVX1 gate1693 ( .A(N6437), .Y(N6905) );
  INVX1 gate1694 ( .A(N6599), .Y(N6908) );
  OR2X1 gate1695 ( .A(N6445), .B(N6194), .Y(N6909) );
  INVX1 gate1696 ( .A(N6606), .Y(N6912) );
  INVX1 gate1697 ( .A(N6609), .Y(N6913) );
  INVX1 gate1698 ( .A(N6619), .Y(N6914) );
  NAND2X1 gate1699 ( .A(N6619), .B(N5734), .Y(N6915) );
  INVX1 gate1700 ( .A(N6445), .Y(N6916) );
  INVX1 gate1701 ( .A(N6622), .Y(N6919) );
  INVX1 gate1702 ( .A(N6634), .Y(N6922) );
  NAND2X1 gate1703 ( .A(N6634), .B(N6067), .Y(N6923) );
  OR2X1 gate1704 ( .A(N6382), .B(N6801), .Y(N6924) );
  OR2X1 gate1705 ( .A(N6386), .B(N6802), .Y(N6925) );
  OR2X1 gate1706 ( .A(N6388), .B(N6803), .Y(N6926) );
  OR2X1 gate1707 ( .A(N6392), .B(N6804), .Y(N6927) );
  INVX1 gate1708 ( .A(N6724), .Y(N6930) );
  NAND2X1 gate1709 ( .A(N6650), .B(N6806), .Y(N6932) );
  NAND2X1 gate1710 ( .A(N6241), .B(N6807), .Y(N6935) );
  NAND2X1 gate1711 ( .A(N6244), .B(N6809), .Y(N6936) );
  NAND2X1 gate1712 ( .A(N6247), .B(N6811), .Y(N6937) );
  NAND2X1 gate1713 ( .A(N6250), .B(N6813), .Y(N6938) );
  NAND2X1 gate1714 ( .A(N6660), .B(N6815), .Y(N6939) );
  NAND2X1 gate1715 ( .A(N6662), .B(N6816), .Y(N6940) );
  NAND2X1 gate1716 ( .A(N6259), .B(N6823), .Y(N6946) );
  NAND2X1 gate1717 ( .A(N6262), .B(N6825), .Y(N6947) );
  NAND2X1 gate1718 ( .A(N6265), .B(N6827), .Y(N6948) );
  NAND2X1 gate1719 ( .A(N6268), .B(N6829), .Y(N6949) );
  NAND2X1 gate1720 ( .A(N5183), .B(N6834), .Y(N6953) );
  NAND2X1 gate1721 ( .A(N5186), .B(N6836), .Y(N6954) );
  NAND2X1 gate1722 ( .A(N5189), .B(N6838), .Y(N6955) );
  NAND2X1 gate1723 ( .A(N5192), .B(N6840), .Y(N6956) );
  NAND2X1 gate1724 ( .A(N6689), .B(N6842), .Y(N6957) );
  NAND2X1 gate1725 ( .A(N6691), .B(N6843), .Y(N6958) );
  NAND2X1 gate1726 ( .A(N6331), .B(N6850), .Y(N6964) );
  NAND2X1 gate1727 ( .A(N6048), .B(N6852), .Y(N6965) );
  NAND2X1 gate1728 ( .A(N6335), .B(N6854), .Y(N6966) );
  NAND2X1 gate1729 ( .A(N6699), .B(N6856), .Y(N6967) );
  NOR2X1 gate1730 ( .A(N6860), .B(N6712), .Y(N6973) );
  NOR2X1 gate1731 ( .A(N6861), .B(N6713), .Y(N6974) );
  NOR2X1 gate1732 ( .A(N6862), .B(N6714), .Y(N6975) );
  NOR2X1 gate1733 ( .A(N6863), .B(N6715), .Y(N6976) );
  INVX1 gate1734 ( .A(N6792), .Y(N6977) );
  INVX1 gate1735 ( .A(N6795), .Y(N6978) );
  OR2X1 gate1736 ( .A(N6879), .B(N6880), .Y(N6979) );
  NAND2X1 gate1737 ( .A(N4608), .B(N6889), .Y(N6987) );
  NAND2X1 gate1738 ( .A(N5177), .B(N6895), .Y(N6990) );
  NAND2X1 gate1739 ( .A(N5217), .B(N6914), .Y(N6999) );
  NAND2X1 gate1740 ( .A(N5377), .B(N6922), .Y(N7002) );
  NAND2X1 gate1741 ( .A(N6873), .B(N6872), .Y(N7003) );
  NAND2X1 gate1742 ( .A(N6875), .B(N6874), .Y(N7006) );
  AND2X1 gate1743_1 ( .A(N6866), .B(N2681), .Y(N7011_1) );
  AND2X1 gate1743 ( .A(N2692), .B(N7011_1), .Y(N7011) );
  AND2X1 gate1744_1 ( .A(N6866), .B(N2756), .Y(N7012_1) );
  AND2X1 gate1744 ( .A(N2767), .B(N7012_1), .Y(N7012) );
  AND2X1 gate1745_1 ( .A(N6866), .B(N2779), .Y(N7013_1) );
  AND2X1 gate1745 ( .A(N2790), .B(N7013_1), .Y(N7013) );
  INVX1 gate1746 ( .A(N6866), .Y(N7015) );
  AND2X1 gate1747_1 ( .A(N6866), .B(N2801), .Y(N7016_1) );
  AND2X1 gate1747 ( .A(N2812), .B(N7016_1), .Y(N7016) );
  NAND2X1 gate1748 ( .A(N6935), .B(N6808), .Y(N7018) );
  NAND2X1 gate1749 ( .A(N6936), .B(N6810), .Y(N7019) );
  NAND2X1 gate1750 ( .A(N6937), .B(N6812), .Y(N7020) );
  NAND2X1 gate1751 ( .A(N6938), .B(N6814), .Y(N7021) );
  INVX1 gate1752 ( .A(N6939), .Y(N7022) );
  INVX1 gate1753 ( .A(N6817), .Y(N7023) );
  NAND2X1 gate1754 ( .A(N6946), .B(N6824), .Y(N7028) );
  NAND2X1 gate1755 ( .A(N6947), .B(N6826), .Y(N7031) );
  NAND2X1 gate1756 ( .A(N6948), .B(N6828), .Y(N7034) );
  NAND2X1 gate1757 ( .A(N6949), .B(N6830), .Y(N7037) );
  AND2X1 gate1758 ( .A(N6817), .B(N6079), .Y(N7040) );
  AND2X1 gate1759 ( .A(N6831), .B(N6675), .Y(N7041) );
  NAND2X1 gate1760 ( .A(N6953), .B(N6835), .Y(N7044) );
  NAND2X1 gate1761 ( .A(N6954), .B(N6837), .Y(N7045) );
  NAND2X1 gate1762 ( .A(N6955), .B(N6839), .Y(N7046) );
  NAND2X1 gate1763 ( .A(N6956), .B(N6841), .Y(N7047) );
  INVX1 gate1764 ( .A(N6957), .Y(N7048) );
  INVX1 gate1765 ( .A(N6844), .Y(N7049) );
  NAND2X1 gate1766 ( .A(N6964), .B(N6851), .Y(N7054) );
  NAND2X1 gate1767 ( .A(N6965), .B(N6853), .Y(N7057) );
  NAND2X1 gate1768 ( .A(N6966), .B(N6855), .Y(N7060) );
  AND2X1 gate1769 ( .A(N6844), .B(N6139), .Y(N7064) );
  AND2X1 gate1770 ( .A(N6857), .B(N6703), .Y(N7065) );
  INVX1 gate1771 ( .A(N6881), .Y(N7072) );
  NAND2X1 gate1772 ( .A(N6881), .B(N5172), .Y(N7073) );
  INVX1 gate1773 ( .A(N6885), .Y(N7074) );
  NAND2X1 gate1774 ( .A(N6885), .B(N5727), .Y(N7075) );
  NAND2X1 gate1775 ( .A(N6890), .B(N6987), .Y(N7076) );
  INVX1 gate1776 ( .A(N6891), .Y(N7079) );
  NAND2X1 gate1777 ( .A(N6896), .B(N6990), .Y(N7080) );
  INVX1 gate1778 ( .A(N6897), .Y(N7083) );
  INVX1 gate1779 ( .A(N6901), .Y(N7084) );
  NAND2X1 gate1780 ( .A(N6901), .B(N5198), .Y(N7085) );
  INVX1 gate1781 ( .A(N6905), .Y(N7086) );
  NAND2X1 gate1782 ( .A(N6905), .B(N5731), .Y(N7087) );
  INVX1 gate1783 ( .A(N6909), .Y(N7088) );
  NAND2X1 gate1784 ( .A(N6909), .B(N6912), .Y(N7089) );
  NAND2X1 gate1785 ( .A(N6915), .B(N6999), .Y(N7090) );
  INVX1 gate1786 ( .A(N6916), .Y(N7093) );
  NAND2X1 gate1787 ( .A(N6974), .B(N6973), .Y(N7094) );
  NAND2X1 gate1788 ( .A(N6976), .B(N6975), .Y(N7097) );
  NAND2X1 gate1789 ( .A(N7002), .B(N6923), .Y(N7101) );
  INVX1 gate1790 ( .A(N6932), .Y(N7105) );
  INVX1 gate1791 ( .A(N6967), .Y(N7110) );
  AND2X1 gate1792_1 ( .A(N6979), .B(N603), .Y(N7114_1) );
  AND2X1 gate1792 ( .A(N1755), .B(N7114_1), .Y(N7114) );
  INVX1 gate1793 ( .A(N7019), .Y(N7115) );
  INVX1 gate1794 ( .A(N7021), .Y(N7116) );
  AND2X1 gate1795 ( .A(N6817), .B(N7018), .Y(N7125) );
  AND2X1 gate1796 ( .A(N6817), .B(N7020), .Y(N7126) );
  AND2X1 gate1797 ( .A(N6817), .B(N7022), .Y(N7127) );
  INVX1 gate1798 ( .A(N7045), .Y(N7130) );
  INVX1 gate1799 ( .A(N7047), .Y(N7131) );
  AND2X1 gate1800 ( .A(N6844), .B(N7044), .Y(N7139) );
  AND2X1 gate1801 ( .A(N6844), .B(N7046), .Y(N7140) );
  AND2X1 gate1802 ( .A(N6844), .B(N7048), .Y(N7141) );
  AND2X1 gate1803_1 ( .A(N6932), .B(N1761), .Y(N7146_1) );
  AND2X1 gate1803 ( .A(N3108), .B(N7146_1), .Y(N7146) );
  AND2X1 gate1804_1 ( .A(N6967), .B(N1777), .Y(N7147_1) );
  AND2X1 gate1804 ( .A(N3130), .B(N7147_1), .Y(N7147) );
  INVX1 gate1805 ( .A(N7003), .Y(N7149) );
  INVX1 gate1806 ( .A(N7006), .Y(N7150) );
  NAND2X1 gate1807 ( .A(N7006), .B(N6876), .Y(N7151) );
  NAND2X1 gate1808 ( .A(N4605), .B(N7072), .Y(N7152) );
  NAND2X1 gate1809 ( .A(N5173), .B(N7074), .Y(N7153) );
  NAND2X1 gate1810 ( .A(N4646), .B(N7084), .Y(N7158) );
  NAND2X1 gate1811 ( .A(N5205), .B(N7086), .Y(N7159) );
  NAND2X1 gate1812 ( .A(N6606), .B(N7088), .Y(N7160) );
  INVX1 gate1813 ( .A(N7037), .Y(N7166) );
  INVX1 gate1814 ( .A(N7034), .Y(N7167) );
  INVX1 gate1815 ( .A(N7031), .Y(N7168) );
  INVX1 gate1816 ( .A(N7028), .Y(N7169) );
  INVX1 gate1817 ( .A(N7060), .Y(N7170) );
  INVX1 gate1818 ( .A(N7057), .Y(N7171) );
  INVX1 gate1819 ( .A(N7054), .Y(N7172) );
  AND2X1 gate1820 ( .A(N7115), .B(N7023), .Y(N7173) );
  AND2X1 gate1821 ( .A(N7116), .B(N7023), .Y(N7174) );
  AND2X1 gate1822 ( .A(N6940), .B(N7023), .Y(N7175) );
  AND2X1 gate1823 ( .A(N5418), .B(N7023), .Y(N7176) );
  INVX1 gate1824 ( .A(N7041), .Y(N7177) );
  AND2X1 gate1825 ( .A(N7130), .B(N7049), .Y(N7178) );
  AND2X1 gate1826 ( .A(N7131), .B(N7049), .Y(N7179) );
  AND2X1 gate1827 ( .A(N6958), .B(N7049), .Y(N7180) );
  AND2X1 gate1828 ( .A(N5573), .B(N7049), .Y(N7181) );
  INVX1 gate1829 ( .A(N7065), .Y(N7182) );
  INVX1 gate1830 ( .A(N7094), .Y(N7183) );
  NAND2X1 gate1831 ( .A(N7094), .B(N6977), .Y(N7184) );
  INVX1 gate1832 ( .A(N7097), .Y(N7185) );
  NAND2X1 gate1833 ( .A(N7097), .B(N6978), .Y(N7186) );
  AND2X1 gate1834_1 ( .A(N7037), .B(N1761), .Y(N7187_1) );
  AND2X1 gate1834 ( .A(N3108), .B(N7187_1), .Y(N7187) );
  AND2X1 gate1835_1 ( .A(N7034), .B(N1761), .Y(N7188_1) );
  AND2X1 gate1835 ( .A(N3108), .B(N7188_1), .Y(N7188) );
  AND2X1 gate1836_1 ( .A(N7031), .B(N1761), .Y(N7189_1) );
  AND2X1 gate1836 ( .A(N3108), .B(N7189_1), .Y(N7189) );
  OR2X1 gate1837_1 ( .A(N4956), .B(N7146), .Y(N7190_1) );
  OR2X1 gate1837 ( .A(N3781), .B(N7190_1), .Y(N7190) );
  AND2X1 gate1838_1 ( .A(N7060), .B(N1777), .Y(N7196_1) );
  AND2X1 gate1838 ( .A(N3130), .B(N7196_1), .Y(N7196) );
  AND2X1 gate1839_1 ( .A(N7057), .B(N1777), .Y(N7197_1) );
  AND2X1 gate1839 ( .A(N3130), .B(N7197_1), .Y(N7197) );
  OR2X1 gate1840_1 ( .A(N4960), .B(N7147), .Y(N7198_1) );
  OR2X1 gate1840 ( .A(N3786), .B(N7198_1), .Y(N7198) );
  NAND2X1 gate1841 ( .A(N7101), .B(N7149), .Y(N7204) );
  INVX1 gate1842 ( .A(N7101), .Y(N7205) );
  NAND2X1 gate1843 ( .A(N6637), .B(N7150), .Y(N7206) );
  AND2X1 gate1844_1 ( .A(N7028), .B(N1793), .Y(N7207_1) );
  AND2X1 gate1844 ( .A(N3158), .B(N7207_1), .Y(N7207) );
  AND2X1 gate1845_1 ( .A(N7054), .B(N1807), .Y(N7208_1) );
  AND2X1 gate1845 ( .A(N3180), .B(N7208_1), .Y(N7208) );
  NAND2X1 gate1846 ( .A(N7073), .B(N7152), .Y(N7209) );
  NAND2X1 gate1847 ( .A(N7075), .B(N7153), .Y(N7212) );
  INVX1 gate1848 ( .A(N7076), .Y(N7215) );
  NAND2X1 gate1849 ( .A(N7076), .B(N7079), .Y(N7216) );
  INVX1 gate1850 ( .A(N7080), .Y(N7217) );
  NAND2X1 gate1851 ( .A(N7080), .B(N7083), .Y(N7218) );
  NAND2X1 gate1852 ( .A(N7085), .B(N7158), .Y(N7219) );
  NAND2X1 gate1853 ( .A(N7087), .B(N7159), .Y(N7222) );
  NAND2X1 gate1854 ( .A(N7089), .B(N7160), .Y(N7225) );
  INVX1 gate1855 ( .A(N7090), .Y(N7228) );
  NAND2X1 gate1856 ( .A(N7090), .B(N7093), .Y(N7229) );
  OR2X1 gate1857 ( .A(N7173), .B(N7125), .Y(N7236) );
  OR2X1 gate1858 ( .A(N7174), .B(N7126), .Y(N7239) );
  OR2X1 gate1859 ( .A(N7175), .B(N7127), .Y(N7242) );
  OR2X1 gate1860 ( .A(N7176), .B(N7040), .Y(N7245) );
  OR2X1 gate1861 ( .A(N7178), .B(N7139), .Y(N7250) );
  OR2X1 gate1862 ( .A(N7179), .B(N7140), .Y(N7257) );
  OR2X1 gate1863 ( .A(N7180), .B(N7141), .Y(N7260) );
  OR2X1 gate1864 ( .A(N7181), .B(N7064), .Y(N7263) );
  NAND2X1 gate1865 ( .A(N6792), .B(N7183), .Y(N7268) );
  NAND2X1 gate1866 ( .A(N6795), .B(N7185), .Y(N7269) );
  OR2X1 gate1867_1 ( .A(N4957), .B(N7187), .Y(N7270_1) );
  OR2X1 gate1867 ( .A(N3782), .B(N7270_1), .Y(N7270) );
  OR2X1 gate1868_1 ( .A(N4958), .B(N7188), .Y(N7276_1) );
  OR2X1 gate1868 ( .A(N3783), .B(N7276_1), .Y(N7276) );
  OR2X1 gate1869_1 ( .A(N4959), .B(N7189), .Y(N7282_1) );
  OR2X1 gate1869 ( .A(N3784), .B(N7282_1), .Y(N7282) );
  OR2X1 gate1870_1 ( .A(N4961), .B(N7196), .Y(N7288_1) );
  OR2X1 gate1870 ( .A(N3787), .B(N7288_1), .Y(N7288) );
  OR2X1 gate1871_1 ( .A(N3998), .B(N7197), .Y(N7294_1) );
  OR2X1 gate1871 ( .A(N3788), .B(N7294_1), .Y(N7294) );
  NAND2X1 gate1872 ( .A(N7003), .B(N7205), .Y(N7300) );
  NAND2X1 gate1873 ( .A(N7206), .B(N7151), .Y(N7301) );
  OR2X1 gate1874_1 ( .A(N4980), .B(N7207), .Y(N7304_1) );
  OR2X1 gate1874 ( .A(N3800), .B(N7304_1), .Y(N7304) );
  OR2X1 gate1875_1 ( .A(N4984), .B(N7208), .Y(N7310_1) );
  OR2X1 gate1875 ( .A(N3805), .B(N7310_1), .Y(N7310) );
  NAND2X1 gate1876 ( .A(N6891), .B(N7215), .Y(N7320) );
  NAND2X1 gate1877 ( .A(N6897), .B(N7217), .Y(N7321) );
  NAND2X1 gate1878 ( .A(N6916), .B(N7228), .Y(N7328) );
  AND2X1 gate1879_1 ( .A(N7190), .B(N1185), .Y(N7338_1) );
  AND2X1 gate1879 ( .A(N2692), .B(N7338_1), .Y(N7338) );
  AND2X1 gate1880_1 ( .A(N7198), .B(N2681), .Y(N7339_1) );
  AND2X1 gate1880 ( .A(N2692), .B(N7339_1), .Y(N7339) );
  AND2X1 gate1881_1 ( .A(N7190), .B(N1247), .Y(N7340_1) );
  AND2X1 gate1881 ( .A(N2767), .B(N7340_1), .Y(N7340) );
  AND2X1 gate1882_1 ( .A(N7198), .B(N2756), .Y(N7341_1) );
  AND2X1 gate1882 ( .A(N2767), .B(N7341_1), .Y(N7341) );
  AND2X1 gate1883_1 ( .A(N7190), .B(N1327), .Y(N7342_1) );
  AND2X1 gate1883 ( .A(N2790), .B(N7342_1), .Y(N7342) );
  AND2X1 gate1884_1 ( .A(N7198), .B(N2779), .Y(N7349_1) );
  AND2X1 gate1884 ( .A(N2790), .B(N7349_1), .Y(N7349) );
  AND2X1 gate1885_1 ( .A(N7198), .B(N2801), .Y(N7357_1) );
  AND2X1 gate1885 ( .A(N2812), .B(N7357_1), .Y(N7357) );
  INVX1 gate1886 ( .A(N7198), .Y(N7363) );
  AND2X1 gate1887_1 ( .A(N7190), .B(N1351), .Y(N7364_1) );
  AND2X1 gate1887 ( .A(N2812), .B(N7364_1), .Y(N7364) );
  INVX1 gate1888 ( .A(N7190), .Y(N7365) );
  NAND2X1 gate1889 ( .A(N7268), .B(N7184), .Y(N7394) );
  NAND2X1 gate1890 ( .A(N7269), .B(N7186), .Y(N7397) );
  NAND2X1 gate1891 ( .A(N7204), .B(N7300), .Y(N7402) );
  INVX1 gate1892 ( .A(N7209), .Y(N7405) );
  NAND2X1 gate1893 ( .A(N7209), .B(N6884), .Y(N7406) );
  INVX1 gate1894 ( .A(N7212), .Y(N7407) );
  NAND2X1 gate1895 ( .A(N7212), .B(N6888), .Y(N7408) );
  NAND2X1 gate1896 ( .A(N7320), .B(N7216), .Y(N7409) );
  NAND2X1 gate1897 ( .A(N7321), .B(N7218), .Y(N7412) );
  INVX1 gate1898 ( .A(N7219), .Y(N7415) );
  NAND2X1 gate1899 ( .A(N7219), .B(N6904), .Y(N7416) );
  INVX1 gate1900 ( .A(N7222), .Y(N7417) );
  NAND2X1 gate1901 ( .A(N7222), .B(N6908), .Y(N7418) );
  INVX1 gate1902 ( .A(N7225), .Y(N7419) );
  NAND2X1 gate1903 ( .A(N7225), .B(N6913), .Y(N7420) );
  NAND2X1 gate1904 ( .A(N7328), .B(N7229), .Y(N7421) );
  INVX1 gate1905 ( .A(N7245), .Y(N7424) );
  INVX1 gate1906 ( .A(N7242), .Y(N7425) );
  INVX1 gate1907 ( .A(N7239), .Y(N7426) );
  INVX1 gate1908 ( .A(N7236), .Y(N7427) );
  INVX1 gate1909 ( .A(N7263), .Y(N7428) );
  INVX1 gate1910 ( .A(N7260), .Y(N7429) );
  INVX1 gate1911 ( .A(N7257), .Y(N7430) );
  INVX1 gate1912 ( .A(N7250), .Y(N7431) );
  INVX1 gate1913 ( .A(N7250), .Y(N7432) );
  AND2X1 gate1914_1 ( .A(N7310), .B(N2653), .Y(N7433_1) );
  AND2X1 gate1914 ( .A(N2664), .B(N7433_1), .Y(N7433) );
  AND2X1 gate1915_1 ( .A(N7304), .B(N1161), .Y(N7434_1) );
  AND2X1 gate1915 ( .A(N2664), .B(N7434_1), .Y(N7434) );
  OR2X1 gate1916_1 ( .A(N7011), .B(N7338), .Y(N7435_1) );
  OR2X1 gate1916_2 ( .A(N3621), .B(N2591), .Y(N7435_2) );
  OR2X1 gate1916 ( .A(N7435_1), .B(N7435_2), .Y(N7435) );
  AND2X1 gate1917_1 ( .A(N7270), .B(N1185), .Y(N7436_1) );
  AND2X1 gate1917 ( .A(N2692), .B(N7436_1), .Y(N7436) );
  AND2X1 gate1918_1 ( .A(N7288), .B(N2681), .Y(N7437_1) );
  AND2X1 gate1918 ( .A(N2692), .B(N7437_1), .Y(N7437) );
  AND2X1 gate1919_1 ( .A(N7276), .B(N1185), .Y(N7438_1) );
  AND2X1 gate1919 ( .A(N2692), .B(N7438_1), .Y(N7438) );
  AND2X1 gate1920_1 ( .A(N7294), .B(N2681), .Y(N7439_1) );
  AND2X1 gate1920 ( .A(N2692), .B(N7439_1), .Y(N7439) );
  AND2X1 gate1921_1 ( .A(N7282), .B(N1185), .Y(N7440_1) );
  AND2X1 gate1921 ( .A(N2692), .B(N7440_1), .Y(N7440) );
  AND2X1 gate1922_1 ( .A(N7310), .B(N2728), .Y(N7441_1) );
  AND2X1 gate1922 ( .A(N2739), .B(N7441_1), .Y(N7441) );
  AND2X1 gate1923_1 ( .A(N7304), .B(N1223), .Y(N7442_1) );
  AND2X1 gate1923 ( .A(N2739), .B(N7442_1), .Y(N7442) );
  OR2X1 gate1924_1 ( .A(N7012), .B(N7340), .Y(N7443_1) );
  OR2X1 gate1924_2 ( .A(N3632), .B(N2600), .Y(N7443_2) );
  OR2X1 gate1924 ( .A(N7443_1), .B(N7443_2), .Y(N7443) );
  AND2X1 gate1925_1 ( .A(N7270), .B(N1247), .Y(N7444_1) );
  AND2X1 gate1925 ( .A(N2767), .B(N7444_1), .Y(N7444) );
  AND2X1 gate1926_1 ( .A(N7288), .B(N2756), .Y(N7445_1) );
  AND2X1 gate1926 ( .A(N2767), .B(N7445_1), .Y(N7445) );
  AND2X1 gate1927_1 ( .A(N7276), .B(N1247), .Y(N7446_1) );
  AND2X1 gate1927 ( .A(N2767), .B(N7446_1), .Y(N7446) );
  AND2X1 gate1928_1 ( .A(N7294), .B(N2756), .Y(N7447_1) );
  AND2X1 gate1928 ( .A(N2767), .B(N7447_1), .Y(N7447) );
  AND2X1 gate1929_1 ( .A(N7282), .B(N1247), .Y(N7448_1) );
  AND2X1 gate1929 ( .A(N2767), .B(N7448_1), .Y(N7448) );
  OR2X1 gate1930_1 ( .A(N7013), .B(N7342), .Y(N7449_1) );
  OR2X1 gate1930_2 ( .A(N3641), .B(N2605), .Y(N7449_2) );
  OR2X1 gate1930 ( .A(N7449_1), .B(N7449_2), .Y(N7449) );
  AND2X1 gate1931_1 ( .A(N7310), .B(N3041), .Y(N7450_1) );
  AND2X1 gate1931 ( .A(N3052), .B(N7450_1), .Y(N7450) );
  AND2X1 gate1932_1 ( .A(N7304), .B(N1697), .Y(N7451_1) );
  AND2X1 gate1932 ( .A(N3052), .B(N7451_1), .Y(N7451) );
  AND2X1 gate1933_1 ( .A(N7294), .B(N2779), .Y(N7452_1) );
  AND2X1 gate1933 ( .A(N2790), .B(N7452_1), .Y(N7452) );
  AND2X1 gate1934_1 ( .A(N7282), .B(N1327), .Y(N7453_1) );
  AND2X1 gate1934 ( .A(N2790), .B(N7453_1), .Y(N7453) );
  AND2X1 gate1935_1 ( .A(N7288), .B(N2779), .Y(N7454_1) );
  AND2X1 gate1935 ( .A(N2790), .B(N7454_1), .Y(N7454) );
  AND2X1 gate1936_1 ( .A(N7276), .B(N1327), .Y(N7455_1) );
  AND2X1 gate1936 ( .A(N2790), .B(N7455_1), .Y(N7455) );
  AND2X1 gate1937_1 ( .A(N7270), .B(N1327), .Y(N7456_1) );
  AND2X1 gate1937 ( .A(N2790), .B(N7456_1), .Y(N7456) );
  AND2X1 gate1938_1 ( .A(N7310), .B(N3075), .Y(N7457_1) );
  AND2X1 gate1938 ( .A(N3086), .B(N7457_1), .Y(N7457) );
  AND2X1 gate1939_1 ( .A(N7304), .B(N1731), .Y(N7458_1) );
  AND2X1 gate1939 ( .A(N3086), .B(N7458_1), .Y(N7458) );
  AND2X1 gate1940_1 ( .A(N7294), .B(N2801), .Y(N7459_1) );
  AND2X1 gate1940 ( .A(N2812), .B(N7459_1), .Y(N7459) );
  AND2X1 gate1941_1 ( .A(N7282), .B(N1351), .Y(N7460_1) );
  AND2X1 gate1941 ( .A(N2812), .B(N7460_1), .Y(N7460) );
  AND2X1 gate1942_1 ( .A(N7288), .B(N2801), .Y(N7461_1) );
  AND2X1 gate1942 ( .A(N2812), .B(N7461_1), .Y(N7461) );
  AND2X1 gate1943_1 ( .A(N7276), .B(N1351), .Y(N7462_1) );
  AND2X1 gate1943 ( .A(N2812), .B(N7462_1), .Y(N7462) );
  AND2X1 gate1944_1 ( .A(N7270), .B(N1351), .Y(N7463_1) );
  AND2X1 gate1944 ( .A(N2812), .B(N7463_1), .Y(N7463) );
  AND2X1 gate1945_1 ( .A(N7250), .B(N603), .Y(N7464_1) );
  AND2X1 gate1945 ( .A(N599), .B(N7464_1), .Y(N7464) );
  INVX1 gate1946 ( .A(N7310), .Y(N7465) );
  INVX1 gate1947 ( .A(N7294), .Y(N7466) );
  INVX1 gate1948 ( .A(N7288), .Y(N7467) );
  INVX1 gate1949 ( .A(N7301), .Y(N7468) );
  OR2X1 gate1950_1 ( .A(N7016), .B(N7364), .Y(N7469_1) );
  OR2X1 gate1950_2 ( .A(N3660), .B(N2626), .Y(N7469_2) );
  OR2X1 gate1950 ( .A(N7469_1), .B(N7469_2), .Y(N7469) );
  INVX1 gate1951 ( .A(N7304), .Y(N7470) );
  INVX1 gate1952 ( .A(N7282), .Y(N7471) );
  INVX1 gate1953 ( .A(N7276), .Y(N7472) );
  INVX1 gate1954 ( .A(N7270), .Y(N7473) );
  BUFX2 gate1955 ( .A(N7394), .Y(N7474) );
  BUFX2 gate1956 ( .A(N7397), .Y(N7476) );
  AND2X1 gate1957 ( .A(N7301), .B(N3068), .Y(N7479) );
  AND2X1 gate1958_1 ( .A(N7245), .B(N1793), .Y(N7481_1) );
  AND2X1 gate1958 ( .A(N3158), .B(N7481_1), .Y(N7481) );
  AND2X1 gate1959_1 ( .A(N7242), .B(N1793), .Y(N7482_1) );
  AND2X1 gate1959 ( .A(N3158), .B(N7482_1), .Y(N7482) );
  AND2X1 gate1960_1 ( .A(N7239), .B(N1793), .Y(N7483_1) );
  AND2X1 gate1960 ( .A(N3158), .B(N7483_1), .Y(N7483) );
  AND2X1 gate1961_1 ( .A(N7236), .B(N1793), .Y(N7484_1) );
  AND2X1 gate1961 ( .A(N3158), .B(N7484_1), .Y(N7484) );
  AND2X1 gate1962_1 ( .A(N7263), .B(N1807), .Y(N7485_1) );
  AND2X1 gate1962 ( .A(N3180), .B(N7485_1), .Y(N7485) );
  AND2X1 gate1963_1 ( .A(N7260), .B(N1807), .Y(N7486_1) );
  AND2X1 gate1963 ( .A(N3180), .B(N7486_1), .Y(N7486) );
  AND2X1 gate1964_1 ( .A(N7257), .B(N1807), .Y(N7487_1) );
  AND2X1 gate1964 ( .A(N3180), .B(N7487_1), .Y(N7487) );
  AND2X1 gate1965_1 ( .A(N7250), .B(N1807), .Y(N7488_1) );
  AND2X1 gate1965 ( .A(N3180), .B(N7488_1), .Y(N7488) );
  NAND2X1 gate1966 ( .A(N6979), .B(N7250), .Y(N7489) );
  NAND2X1 gate1967 ( .A(N6516), .B(N7405), .Y(N7492) );
  NAND2X1 gate1968 ( .A(N6526), .B(N7407), .Y(N7493) );
  NAND2X1 gate1969 ( .A(N6592), .B(N7415), .Y(N7498) );
  NAND2X1 gate1970 ( .A(N6599), .B(N7417), .Y(N7499) );
  NAND2X1 gate1971 ( .A(N6609), .B(N7419), .Y(N7500) );
  AND2X1 gate1972_1 ( .A(N7105), .B(N7166), .Y(N7503_1) );
  AND2X1 gate1972_2 ( .A(N7167), .B(N7168), .Y(N7503_2) );
  AND2X1 gate1972_3 ( .A(N7169), .B(N7424), .Y(N7503_3) );
  AND2X1 gate1972_4 ( .A(N7425), .B(N7426), .Y(N7503_4) );
  AND2X1 gate1972_5 ( .A(N7427), .B(N7503_1), .Y(N7503_5) );
  AND2X1 gate1972_6 ( .A(N7503_2), .B(N7503_3), .Y(N7503_6) );
  AND2X1 gate1972_7 ( .A(N7503_4), .B(N7503_5), .Y(N7503_7) );
  AND2X1 gate1972 ( .A(N7503_6), .B(N7503_7), .Y(N7503) );
  AND2X1 gate1973_1 ( .A(N6640), .B(N7110), .Y(N7504_1) );
  AND2X1 gate1973_2 ( .A(N7170), .B(N7171), .Y(N7504_2) );
  AND2X1 gate1973_3 ( .A(N7172), .B(N7428), .Y(N7504_3) );
  AND2X1 gate1973_4 ( .A(N7429), .B(N7430), .Y(N7504_4) );
  AND2X1 gate1973_5 ( .A(N7431), .B(N7504_1), .Y(N7504_5) );
  AND2X1 gate1973_6 ( .A(N7504_2), .B(N7504_3), .Y(N7504_6) );
  AND2X1 gate1973_7 ( .A(N7504_4), .B(N7504_5), .Y(N7504_7) );
  AND2X1 gate1973 ( .A(N7504_6), .B(N7504_7), .Y(N7504) );
  OR2X1 gate1974_1 ( .A(N7433), .B(N7434), .Y(N7505_1) );
  OR2X1 gate1974_2 ( .A(N3616), .B(N2585), .Y(N7505_2) );
  OR2X1 gate1974 ( .A(N7505_1), .B(N7505_2), .Y(N7505) );
  AND2X1 gate1975 ( .A(N7435), .B(N2675), .Y(N7506) );
  OR2X1 gate1976_1 ( .A(N7339), .B(N7436), .Y(N7507_1) );
  OR2X1 gate1976_2 ( .A(N3622), .B(N2592), .Y(N7507_2) );
  OR2X1 gate1976 ( .A(N7507_1), .B(N7507_2), .Y(N7507) );
  OR2X1 gate1977_1 ( .A(N7437), .B(N7438), .Y(N7508_1) );
  OR2X1 gate1977_2 ( .A(N3623), .B(N2593), .Y(N7508_2) );
  OR2X1 gate1977 ( .A(N7508_1), .B(N7508_2), .Y(N7508) );
  OR2X1 gate1978_1 ( .A(N7439), .B(N7440), .Y(N7509_1) );
  OR2X1 gate1978_2 ( .A(N3624), .B(N2594), .Y(N7509_2) );
  OR2X1 gate1978 ( .A(N7509_1), .B(N7509_2), .Y(N7509) );
  OR2X1 gate1979_1 ( .A(N7441), .B(N7442), .Y(N7510_1) );
  OR2X1 gate1979_2 ( .A(N3627), .B(N2595), .Y(N7510_2) );
  OR2X1 gate1979 ( .A(N7510_1), .B(N7510_2), .Y(N7510) );
  AND2X1 gate1980 ( .A(N7443), .B(N2750), .Y(N7511) );
  OR2X1 gate1981_1 ( .A(N7341), .B(N7444), .Y(N7512_1) );
  OR2X1 gate1981_2 ( .A(N3633), .B(N2601), .Y(N7512_2) );
  OR2X1 gate1981 ( .A(N7512_1), .B(N7512_2), .Y(N7512) );
  OR2X1 gate1982_1 ( .A(N7445), .B(N7446), .Y(N7513_1) );
  OR2X1 gate1982_2 ( .A(N3634), .B(N2602), .Y(N7513_2) );
  OR2X1 gate1982 ( .A(N7513_1), .B(N7513_2), .Y(N7513) );
  OR2X1 gate1983_1 ( .A(N7447), .B(N7448), .Y(N7514_1) );
  OR2X1 gate1983_2 ( .A(N3635), .B(N2603), .Y(N7514_2) );
  OR2X1 gate1983 ( .A(N7514_1), .B(N7514_2), .Y(N7514) );
  OR2X1 gate1984_1 ( .A(N7450), .B(N7451), .Y(N7515_1) );
  OR2X1 gate1984_2 ( .A(N3646), .B(N2610), .Y(N7515_2) );
  OR2X1 gate1984 ( .A(N7515_1), .B(N7515_2), .Y(N7515) );
  OR2X1 gate1985_1 ( .A(N7452), .B(N7453), .Y(N7516_1) );
  OR2X1 gate1985_2 ( .A(N3647), .B(N2611), .Y(N7516_2) );
  OR2X1 gate1985 ( .A(N7516_1), .B(N7516_2), .Y(N7516) );
  OR2X1 gate1986_1 ( .A(N7454), .B(N7455), .Y(N7517_1) );
  OR2X1 gate1986_2 ( .A(N3648), .B(N2612), .Y(N7517_2) );
  OR2X1 gate1986 ( .A(N7517_1), .B(N7517_2), .Y(N7517) );
  OR2X1 gate1987_1 ( .A(N7349), .B(N7456), .Y(N7518_1) );
  OR2X1 gate1987_2 ( .A(N3649), .B(N2613), .Y(N7518_2) );
  OR2X1 gate1987 ( .A(N7518_1), .B(N7518_2), .Y(N7518) );
  OR2X1 gate1988_1 ( .A(N7457), .B(N7458), .Y(N7519_1) );
  OR2X1 gate1988_2 ( .A(N3654), .B(N2618), .Y(N7519_2) );
  OR2X1 gate1988 ( .A(N7519_1), .B(N7519_2), .Y(N7519) );
  OR2X1 gate1989_1 ( .A(N7459), .B(N7460), .Y(N7520_1) );
  OR2X1 gate1989_2 ( .A(N3655), .B(N2619), .Y(N7520_2) );
  OR2X1 gate1989 ( .A(N7520_1), .B(N7520_2), .Y(N7520) );
  OR2X1 gate1990_1 ( .A(N7461), .B(N7462), .Y(N7521_1) );
  OR2X1 gate1990_2 ( .A(N3656), .B(N2620), .Y(N7521_2) );
  OR2X1 gate1990 ( .A(N7521_1), .B(N7521_2), .Y(N7521) );
  OR2X1 gate1991_1 ( .A(N7357), .B(N7463), .Y(N7522_1) );
  OR2X1 gate1991_2 ( .A(N3657), .B(N2621), .Y(N7522_2) );
  OR2X1 gate1991 ( .A(N7522_1), .B(N7522_2), .Y(N7522) );
  OR2X1 gate1992_1 ( .A(N4741), .B(N7114), .Y(N7525_1) );
  OR2X1 gate1992_2 ( .A(N2624), .B(N7464), .Y(N7525_2) );
  OR2X1 gate1992 ( .A(N7525_1), .B(N7525_2), .Y(N7525) );
  AND2X1 gate1993_1 ( .A(N7468), .B(N3119), .Y(N7526_1) );
  AND2X1 gate1993 ( .A(N3130), .B(N7526_1), .Y(N7526) );
  INVX1 gate1994 ( .A(N7394), .Y(N7527) );
  INVX1 gate1995 ( .A(N7397), .Y(N7528) );
  INVX1 gate1996 ( .A(N7402), .Y(N7529) );
  AND2X1 gate1997 ( .A(N7402), .B(N3068), .Y(N7530) );
  OR2X1 gate1998_1 ( .A(N4981), .B(N7481), .Y(N7531_1) );
  OR2X1 gate1998 ( .A(N3801), .B(N7531_1), .Y(N7531) );
  OR2X1 gate1999_1 ( .A(N4982), .B(N7482), .Y(N7537_1) );
  OR2X1 gate1999 ( .A(N3802), .B(N7537_1), .Y(N7537) );
  OR2X1 gate2000_1 ( .A(N4983), .B(N7483), .Y(N7543_1) );
  OR2X1 gate2000 ( .A(N3803), .B(N7543_1), .Y(N7543) );
  OR2X1 gate2001_1 ( .A(N5165), .B(N7484), .Y(N7549_1) );
  OR2X1 gate2001 ( .A(N3804), .B(N7549_1), .Y(N7549) );
  OR2X1 gate2002_1 ( .A(N4985), .B(N7485), .Y(N7555_1) );
  OR2X1 gate2002 ( .A(N3806), .B(N7555_1), .Y(N7555) );
  OR2X1 gate2003_1 ( .A(N4986), .B(N7486), .Y(N7561_1) );
  OR2X1 gate2003 ( .A(N3807), .B(N7561_1), .Y(N7561) );
  OR2X1 gate2004_1 ( .A(N4547), .B(N7487), .Y(N7567_1) );
  OR2X1 gate2004 ( .A(N3808), .B(N7567_1), .Y(N7567) );
  OR2X1 gate2005_1 ( .A(N4987), .B(N7488), .Y(N7573_1) );
  OR2X1 gate2005 ( .A(N3809), .B(N7573_1), .Y(N7573) );
  NAND2X1 gate2006 ( .A(N7492), .B(N7406), .Y(N7579) );
  NAND2X1 gate2007 ( .A(N7493), .B(N7408), .Y(N7582) );
  INVX1 gate2008 ( .A(N7409), .Y(N7585) );
  NAND2X1 gate2009 ( .A(N7409), .B(N6894), .Y(N7586) );
  INVX1 gate2010 ( .A(N7412), .Y(N7587) );
  NAND2X1 gate2011 ( .A(N7412), .B(N6900), .Y(N7588) );
  NAND2X1 gate2012 ( .A(N7498), .B(N7416), .Y(N7589) );
  NAND2X1 gate2013 ( .A(N7499), .B(N7418), .Y(N7592) );
  NAND2X1 gate2014 ( .A(N7500), .B(N7420), .Y(N7595) );
  INVX1 gate2015 ( .A(N7421), .Y(N7598) );
  NAND2X1 gate2016 ( .A(N7421), .B(N6919), .Y(N7599) );
  AND2X1 gate2017 ( .A(N7505), .B(N2647), .Y(N7600) );
  AND2X1 gate2018 ( .A(N7507), .B(N2675), .Y(N7601) );
  AND2X1 gate2019 ( .A(N7508), .B(N2675), .Y(N7602) );
  AND2X1 gate2020 ( .A(N7509), .B(N2675), .Y(N7603) );
  AND2X1 gate2021 ( .A(N7510), .B(N2722), .Y(N7604) );
  AND2X1 gate2022 ( .A(N7512), .B(N2750), .Y(N7605) );
  AND2X1 gate2023 ( .A(N7513), .B(N2750), .Y(N7606) );
  AND2X1 gate2024 ( .A(N7514), .B(N2750), .Y(N7607) );
  AND2X1 gate2025 ( .A(N6979), .B(N7489), .Y(N7624) );
  AND2X1 gate2026 ( .A(N7489), .B(N7250), .Y(N7625) );
  AND2X1 gate2027 ( .A(N1149), .B(N7525), .Y(N7626) );
  AND2X1 gate2028_1 ( .A(N562), .B(N7527), .Y(N7631_1) );
  AND2X1 gate2028_2 ( .A(N7528), .B(N6805), .Y(N7631_2) );
  AND2X1 gate2028_3 ( .A(N6930), .B(N7631_1), .Y(N7631_3) );
  AND2X1 gate2028 ( .A(N7631_2), .B(N7631_3), .Y(N7631) );
  AND2X1 gate2029_1 ( .A(N7529), .B(N3097), .Y(N7636_1) );
  AND2X1 gate2029 ( .A(N3108), .B(N7636_1), .Y(N7636) );
  NAND2X1 gate2030 ( .A(N6539), .B(N7585), .Y(N7657) );
  NAND2X1 gate2031 ( .A(N6556), .B(N7587), .Y(N7658) );
  NAND2X1 gate2032 ( .A(N6622), .B(N7598), .Y(N7665) );
  AND2X1 gate2033_1 ( .A(N7555), .B(N2653), .Y(N7666_1) );
  AND2X1 gate2033 ( .A(N2664), .B(N7666_1), .Y(N7666) );
  AND2X1 gate2034_1 ( .A(N7531), .B(N1161), .Y(N7667_1) );
  AND2X1 gate2034 ( .A(N2664), .B(N7667_1), .Y(N7667) );
  AND2X1 gate2035_1 ( .A(N7561), .B(N2653), .Y(N7668_1) );
  AND2X1 gate2035 ( .A(N2664), .B(N7668_1), .Y(N7668) );
  AND2X1 gate2036_1 ( .A(N7537), .B(N1161), .Y(N7669_1) );
  AND2X1 gate2036 ( .A(N2664), .B(N7669_1), .Y(N7669) );
  AND2X1 gate2037_1 ( .A(N7567), .B(N2653), .Y(N7670_1) );
  AND2X1 gate2037 ( .A(N2664), .B(N7670_1), .Y(N7670) );
  AND2X1 gate2038_1 ( .A(N7543), .B(N1161), .Y(N7671_1) );
  AND2X1 gate2038 ( .A(N2664), .B(N7671_1), .Y(N7671) );
  AND2X1 gate2039_1 ( .A(N7573), .B(N2653), .Y(N7672_1) );
  AND2X1 gate2039 ( .A(N2664), .B(N7672_1), .Y(N7672) );
  AND2X1 gate2040_1 ( .A(N7549), .B(N1161), .Y(N7673_1) );
  AND2X1 gate2040 ( .A(N2664), .B(N7673_1), .Y(N7673) );
  AND2X1 gate2041_1 ( .A(N7555), .B(N2728), .Y(N7674_1) );
  AND2X1 gate2041 ( .A(N2739), .B(N7674_1), .Y(N7674) );
  AND2X1 gate2042_1 ( .A(N7531), .B(N1223), .Y(N7675_1) );
  AND2X1 gate2042 ( .A(N2739), .B(N7675_1), .Y(N7675) );
  AND2X1 gate2043_1 ( .A(N7561), .B(N2728), .Y(N7676_1) );
  AND2X1 gate2043 ( .A(N2739), .B(N7676_1), .Y(N7676) );
  AND2X1 gate2044_1 ( .A(N7537), .B(N1223), .Y(N7677_1) );
  AND2X1 gate2044 ( .A(N2739), .B(N7677_1), .Y(N7677) );
  AND2X1 gate2045_1 ( .A(N7567), .B(N2728), .Y(N7678_1) );
  AND2X1 gate2045 ( .A(N2739), .B(N7678_1), .Y(N7678) );
  AND2X1 gate2046_1 ( .A(N7543), .B(N1223), .Y(N7679_1) );
  AND2X1 gate2046 ( .A(N2739), .B(N7679_1), .Y(N7679) );
  AND2X1 gate2047_1 ( .A(N7573), .B(N2728), .Y(N7680_1) );
  AND2X1 gate2047 ( .A(N2739), .B(N7680_1), .Y(N7680) );
  AND2X1 gate2048_1 ( .A(N7549), .B(N1223), .Y(N7681_1) );
  AND2X1 gate2048 ( .A(N2739), .B(N7681_1), .Y(N7681) );
  AND2X1 gate2049_1 ( .A(N7573), .B(N3075), .Y(N7682_1) );
  AND2X1 gate2049 ( .A(N3086), .B(N7682_1), .Y(N7682) );
  AND2X1 gate2050_1 ( .A(N7549), .B(N1731), .Y(N7683_1) );
  AND2X1 gate2050 ( .A(N3086), .B(N7683_1), .Y(N7683) );
  AND2X1 gate2051_1 ( .A(N7573), .B(N3041), .Y(N7684_1) );
  AND2X1 gate2051 ( .A(N3052), .B(N7684_1), .Y(N7684) );
  AND2X1 gate2052_1 ( .A(N7549), .B(N1697), .Y(N7685_1) );
  AND2X1 gate2052 ( .A(N3052), .B(N7685_1), .Y(N7685) );
  AND2X1 gate2053_1 ( .A(N7567), .B(N3041), .Y(N7686_1) );
  AND2X1 gate2053 ( .A(N3052), .B(N7686_1), .Y(N7686) );
  AND2X1 gate2054_1 ( .A(N7543), .B(N1697), .Y(N7687_1) );
  AND2X1 gate2054 ( .A(N3052), .B(N7687_1), .Y(N7687) );
  AND2X1 gate2055_1 ( .A(N7561), .B(N3041), .Y(N7688_1) );
  AND2X1 gate2055 ( .A(N3052), .B(N7688_1), .Y(N7688) );
  AND2X1 gate2056_1 ( .A(N7537), .B(N1697), .Y(N7689_1) );
  AND2X1 gate2056 ( .A(N3052), .B(N7689_1), .Y(N7689) );
  AND2X1 gate2057_1 ( .A(N7555), .B(N3041), .Y(N7690_1) );
  AND2X1 gate2057 ( .A(N3052), .B(N7690_1), .Y(N7690) );
  AND2X1 gate2058_1 ( .A(N7531), .B(N1697), .Y(N7691_1) );
  AND2X1 gate2058 ( .A(N3052), .B(N7691_1), .Y(N7691) );
  AND2X1 gate2059_1 ( .A(N7567), .B(N3075), .Y(N7692_1) );
  AND2X1 gate2059 ( .A(N3086), .B(N7692_1), .Y(N7692) );
  AND2X1 gate2060_1 ( .A(N7543), .B(N1731), .Y(N7693_1) );
  AND2X1 gate2060 ( .A(N3086), .B(N7693_1), .Y(N7693) );
  AND2X1 gate2061_1 ( .A(N7561), .B(N3075), .Y(N7694_1) );
  AND2X1 gate2061 ( .A(N3086), .B(N7694_1), .Y(N7694) );
  AND2X1 gate2062_1 ( .A(N7537), .B(N1731), .Y(N7695_1) );
  AND2X1 gate2062 ( .A(N3086), .B(N7695_1), .Y(N7695) );
  AND2X1 gate2063_1 ( .A(N7555), .B(N3075), .Y(N7696_1) );
  AND2X1 gate2063 ( .A(N3086), .B(N7696_1), .Y(N7696) );
  AND2X1 gate2064_1 ( .A(N7531), .B(N1731), .Y(N7697_1) );
  AND2X1 gate2064 ( .A(N3086), .B(N7697_1), .Y(N7697) );
  OR2X1 gate2065 ( .A(N7624), .B(N7625), .Y(N7698) );
  INVX1 gate2066 ( .A(N7573), .Y(N7699) );
  INVX1 gate2067 ( .A(N7567), .Y(N7700) );
  INVX1 gate2068 ( .A(N7561), .Y(N7701) );
  INVX1 gate2069 ( .A(N7555), .Y(N7702) );
  AND2X1 gate2070_1 ( .A(N1156), .B(N7631), .Y(N7703_1) );
  AND2X1 gate2070 ( .A(N245), .B(N7703_1), .Y(N7703) );
  INVX1 gate2071 ( .A(N7549), .Y(N7704) );
  INVX1 gate2072 ( .A(N7543), .Y(N7705) );
  INVX1 gate2073 ( .A(N7537), .Y(N7706) );
  INVX1 gate2074 ( .A(N7531), .Y(N7707) );
  INVX1 gate2075 ( .A(N7579), .Y(N7708) );
  NAND2X1 gate2076 ( .A(N7579), .B(N6739), .Y(N7709) );
  INVX1 gate2077 ( .A(N7582), .Y(N7710) );
  NAND2X1 gate2078 ( .A(N7582), .B(N6744), .Y(N7711) );
  NAND2X1 gate2079 ( .A(N7657), .B(N7586), .Y(N7712) );
  NAND2X1 gate2080 ( .A(N7658), .B(N7588), .Y(N7715) );
  INVX1 gate2081 ( .A(N7589), .Y(N7718) );
  NAND2X1 gate2082 ( .A(N7589), .B(N6772), .Y(N7719) );
  INVX1 gate2083 ( .A(N7592), .Y(N7720) );
  NAND2X1 gate2084 ( .A(N7592), .B(N6776), .Y(N7721) );
  INVX1 gate2085 ( .A(N7595), .Y(N7722) );
  NAND2X1 gate2086 ( .A(N7595), .B(N5733), .Y(N7723) );
  NAND2X1 gate2087 ( .A(N7665), .B(N7599), .Y(N7724) );
  OR2X1 gate2088_1 ( .A(N7666), .B(N7667), .Y(N7727_1) );
  OR2X1 gate2088_2 ( .A(N3617), .B(N2586), .Y(N7727_2) );
  OR2X1 gate2088 ( .A(N7727_1), .B(N7727_2), .Y(N7727) );
  OR2X1 gate2089_1 ( .A(N7668), .B(N7669), .Y(N7728_1) );
  OR2X1 gate2089_2 ( .A(N3618), .B(N2587), .Y(N7728_2) );
  OR2X1 gate2089 ( .A(N7728_1), .B(N7728_2), .Y(N7728) );
  OR2X1 gate2090_1 ( .A(N7670), .B(N7671), .Y(N7729_1) );
  OR2X1 gate2090_2 ( .A(N3619), .B(N2588), .Y(N7729_2) );
  OR2X1 gate2090 ( .A(N7729_1), .B(N7729_2), .Y(N7729) );
  OR2X1 gate2091_1 ( .A(N7672), .B(N7673), .Y(N7730_1) );
  OR2X1 gate2091_2 ( .A(N3620), .B(N2589), .Y(N7730_2) );
  OR2X1 gate2091 ( .A(N7730_1), .B(N7730_2), .Y(N7730) );
  OR2X1 gate2092_1 ( .A(N7674), .B(N7675), .Y(N7731_1) );
  OR2X1 gate2092_2 ( .A(N3628), .B(N2596), .Y(N7731_2) );
  OR2X1 gate2092 ( .A(N7731_1), .B(N7731_2), .Y(N7731) );
  OR2X1 gate2093_1 ( .A(N7676), .B(N7677), .Y(N7732_1) );
  OR2X1 gate2093_2 ( .A(N3629), .B(N2597), .Y(N7732_2) );
  OR2X1 gate2093 ( .A(N7732_1), .B(N7732_2), .Y(N7732) );
  OR2X1 gate2094_1 ( .A(N7678), .B(N7679), .Y(N7733_1) );
  OR2X1 gate2094_2 ( .A(N3630), .B(N2598), .Y(N7733_2) );
  OR2X1 gate2094 ( .A(N7733_1), .B(N7733_2), .Y(N7733) );
  OR2X1 gate2095_1 ( .A(N7680), .B(N7681), .Y(N7734_1) );
  OR2X1 gate2095_2 ( .A(N3631), .B(N2599), .Y(N7734_2) );
  OR2X1 gate2095 ( .A(N7734_1), .B(N7734_2), .Y(N7734) );
  OR2X1 gate2096_1 ( .A(N7682), .B(N7683), .Y(N7735_1) );
  OR2X1 gate2096_2 ( .A(N3638), .B(N2604), .Y(N7735_2) );
  OR2X1 gate2096 ( .A(N7735_1), .B(N7735_2), .Y(N7735) );
  OR2X1 gate2097_1 ( .A(N7684), .B(N7685), .Y(N7736_1) );
  OR2X1 gate2097_2 ( .A(N3642), .B(N2606), .Y(N7736_2) );
  OR2X1 gate2097 ( .A(N7736_1), .B(N7736_2), .Y(N7736) );
  OR2X1 gate2098_1 ( .A(N7686), .B(N7687), .Y(N7737_1) );
  OR2X1 gate2098_2 ( .A(N3643), .B(N2607), .Y(N7737_2) );
  OR2X1 gate2098 ( .A(N7737_1), .B(N7737_2), .Y(N7737) );
  OR2X1 gate2099_1 ( .A(N7688), .B(N7689), .Y(N7738_1) );
  OR2X1 gate2099_2 ( .A(N3644), .B(N2608), .Y(N7738_2) );
  OR2X1 gate2099 ( .A(N7738_1), .B(N7738_2), .Y(N7738) );
  OR2X1 gate2100_1 ( .A(N7690), .B(N7691), .Y(N7739_1) );
  OR2X1 gate2100_2 ( .A(N3645), .B(N2609), .Y(N7739_2) );
  OR2X1 gate2100 ( .A(N7739_1), .B(N7739_2), .Y(N7739) );
  OR2X1 gate2101_1 ( .A(N7692), .B(N7693), .Y(N7740_1) );
  OR2X1 gate2101_2 ( .A(N3651), .B(N2615), .Y(N7740_2) );
  OR2X1 gate2101 ( .A(N7740_1), .B(N7740_2), .Y(N7740) );
  OR2X1 gate2102_1 ( .A(N7694), .B(N7695), .Y(N7741_1) );
  OR2X1 gate2102_2 ( .A(N3652), .B(N2616), .Y(N7741_2) );
  OR2X1 gate2102 ( .A(N7741_1), .B(N7741_2), .Y(N7741) );
  OR2X1 gate2103_1 ( .A(N7696), .B(N7697), .Y(N7742_1) );
  OR2X1 gate2103_2 ( .A(N3653), .B(N2617), .Y(N7742_2) );
  OR2X1 gate2103 ( .A(N7742_1), .B(N7742_2), .Y(N7742) );
  NAND2X1 gate2104 ( .A(N6271), .B(N7708), .Y(N7743) );
  NAND2X1 gate2105 ( .A(N6283), .B(N7710), .Y(N7744) );
  NAND2X1 gate2106 ( .A(N6341), .B(N7718), .Y(N7749) );
  NAND2X1 gate2107 ( .A(N6347), .B(N7720), .Y(N7750) );
  NAND2X1 gate2108 ( .A(N5214), .B(N7722), .Y(N7751) );
  AND2X1 gate2109 ( .A(N7727), .B(N2647), .Y(N7754) );
  AND2X1 gate2110 ( .A(N7728), .B(N2647), .Y(N7755) );
  AND2X1 gate2111 ( .A(N7729), .B(N2647), .Y(N7756) );
  AND2X1 gate2112 ( .A(N7730), .B(N2647), .Y(N7757) );
  AND2X1 gate2113 ( .A(N7731), .B(N2722), .Y(N7758) );
  AND2X1 gate2114 ( .A(N7732), .B(N2722), .Y(N7759) );
  AND2X1 gate2115 ( .A(N7733), .B(N2722), .Y(N7760) );
  AND2X1 gate2116 ( .A(N7734), .B(N2722), .Y(N7761) );
  NAND2X1 gate2117 ( .A(N7743), .B(N7709), .Y(N7762) );
  NAND2X1 gate2118 ( .A(N7744), .B(N7711), .Y(N7765) );
  INVX1 gate2119 ( .A(N7712), .Y(N7768) );
  NAND2X1 gate2120 ( .A(N7712), .B(N6751), .Y(N7769) );
  INVX1 gate2121 ( .A(N7715), .Y(N7770) );
  NAND2X1 gate2122 ( .A(N7715), .B(N6760), .Y(N7771) );
  NAND2X1 gate2123 ( .A(N7749), .B(N7719), .Y(N7772) );
  NAND2X1 gate2124 ( .A(N7750), .B(N7721), .Y(N7775) );
  NAND2X1 gate2125 ( .A(N7751), .B(N7723), .Y(N7778) );
  INVX1 gate2126 ( .A(N7724), .Y(N7781) );
  NAND2X1 gate2127 ( .A(N7724), .B(N5735), .Y(N7782) );
  NAND2X1 gate2128 ( .A(N6295), .B(N7768), .Y(N7787) );
  NAND2X1 gate2129 ( .A(N6313), .B(N7770), .Y(N7788) );
  NAND2X1 gate2130 ( .A(N5220), .B(N7781), .Y(N7795) );
  INVX1 gate2131 ( .A(N7762), .Y(N7796) );
  NAND2X1 gate2132 ( .A(N7762), .B(N6740), .Y(N7797) );
  INVX1 gate2133 ( .A(N7765), .Y(N7798) );
  NAND2X1 gate2134 ( .A(N7765), .B(N6745), .Y(N7799) );
  NAND2X1 gate2135 ( .A(N7787), .B(N7769), .Y(N7800) );
  NAND2X1 gate2136 ( .A(N7788), .B(N7771), .Y(N7803) );
  INVX1 gate2137 ( .A(N7772), .Y(N7806) );
  NAND2X1 gate2138 ( .A(N7772), .B(N6773), .Y(N7807) );
  INVX1 gate2139 ( .A(N7775), .Y(N7808) );
  NAND2X1 gate2140 ( .A(N7775), .B(N6777), .Y(N7809) );
  INVX1 gate2141 ( .A(N7778), .Y(N7810) );
  NAND2X1 gate2142 ( .A(N7778), .B(N6782), .Y(N7811) );
  NAND2X1 gate2143 ( .A(N7795), .B(N7782), .Y(N7812) );
  NAND2X1 gate2144 ( .A(N6274), .B(N7796), .Y(N7815) );
  NAND2X1 gate2145 ( .A(N6286), .B(N7798), .Y(N7816) );
  NAND2X1 gate2146 ( .A(N6344), .B(N7806), .Y(N7821) );
  NAND2X1 gate2147 ( .A(N6350), .B(N7808), .Y(N7822) );
  NAND2X1 gate2148 ( .A(N6353), .B(N7810), .Y(N7823) );
  NAND2X1 gate2149 ( .A(N7815), .B(N7797), .Y(N7826) );
  NAND2X1 gate2150 ( .A(N7816), .B(N7799), .Y(N7829) );
  INVX1 gate2151 ( .A(N7800), .Y(N7832) );
  NAND2X1 gate2152 ( .A(N7800), .B(N6752), .Y(N7833) );
  INVX1 gate2153 ( .A(N7803), .Y(N7834) );
  NAND2X1 gate2154 ( .A(N7803), .B(N6761), .Y(N7835) );
  NAND2X1 gate2155 ( .A(N7821), .B(N7807), .Y(N7836) );
  NAND2X1 gate2156 ( .A(N7822), .B(N7809), .Y(N7839) );
  NAND2X1 gate2157 ( .A(N7823), .B(N7811), .Y(N7842) );
  INVX1 gate2158 ( .A(N7812), .Y(N7845) );
  NAND2X1 gate2159 ( .A(N7812), .B(N6790), .Y(N7846) );
  NAND2X1 gate2160 ( .A(N6298), .B(N7832), .Y(N7851) );
  NAND2X1 gate2161 ( .A(N6316), .B(N7834), .Y(N7852) );
  NAND2X1 gate2162 ( .A(N6364), .B(N7845), .Y(N7859) );
  INVX1 gate2163 ( .A(N7826), .Y(N7860) );
  NAND2X1 gate2164 ( .A(N7826), .B(N6741), .Y(N7861) );
  INVX1 gate2165 ( .A(N7829), .Y(N7862) );
  NAND2X1 gate2166 ( .A(N7829), .B(N6746), .Y(N7863) );
  NAND2X1 gate2167 ( .A(N7851), .B(N7833), .Y(N7864) );
  NAND2X1 gate2168 ( .A(N7852), .B(N7835), .Y(N7867) );
  INVX1 gate2169 ( .A(N7836), .Y(N7870) );
  NAND2X1 gate2170 ( .A(N7836), .B(N5730), .Y(N7871) );
  INVX1 gate2171 ( .A(N7839), .Y(N7872) );
  NAND2X1 gate2172 ( .A(N7839), .B(N5732), .Y(N7873) );
  INVX1 gate2173 ( .A(N7842), .Y(N7874) );
  NAND2X1 gate2174 ( .A(N7842), .B(N6783), .Y(N7875) );
  NAND2X1 gate2175 ( .A(N7859), .B(N7846), .Y(N7876) );
  NAND2X1 gate2176 ( .A(N6277), .B(N7860), .Y(N7879) );
  NAND2X1 gate2177 ( .A(N6289), .B(N7862), .Y(N7880) );
  NAND2X1 gate2178 ( .A(N5199), .B(N7870), .Y(N7885) );
  NAND2X1 gate2179 ( .A(N5208), .B(N7872), .Y(N7886) );
  NAND2X1 gate2180 ( .A(N6356), .B(N7874), .Y(N7887) );
  NAND2X1 gate2181 ( .A(N7879), .B(N7861), .Y(N7890) );
  NAND2X1 gate2182 ( .A(N7880), .B(N7863), .Y(N7893) );
  INVX1 gate2183 ( .A(N7864), .Y(N7896) );
  NAND2X1 gate2184 ( .A(N7864), .B(N6753), .Y(N7897) );
  INVX1 gate2185 ( .A(N7867), .Y(N7898) );
  NAND2X1 gate2186 ( .A(N7867), .B(N6762), .Y(N7899) );
  NAND2X1 gate2187 ( .A(N7885), .B(N7871), .Y(N7900) );
  NAND2X1 gate2188 ( .A(N7886), .B(N7873), .Y(N7903) );
  NAND2X1 gate2189 ( .A(N7887), .B(N7875), .Y(N7906) );
  INVX1 gate2190 ( .A(N7876), .Y(N7909) );
  NAND2X1 gate2191 ( .A(N7876), .B(N6791), .Y(N7910) );
  NAND2X1 gate2192 ( .A(N6301), .B(N7896), .Y(N7917) );
  NAND2X1 gate2193 ( .A(N6319), .B(N7898), .Y(N7918) );
  NAND2X1 gate2194 ( .A(N6367), .B(N7909), .Y(N7923) );
  INVX1 gate2195 ( .A(N7890), .Y(N7924) );
  NAND2X1 gate2196 ( .A(N7890), .B(N6680), .Y(N7925) );
  INVX1 gate2197 ( .A(N7893), .Y(N7926) );
  NAND2X1 gate2198 ( .A(N7893), .B(N6681), .Y(N7927) );
  INVX1 gate2199 ( .A(N7900), .Y(N7928) );
  NAND2X1 gate2200 ( .A(N7900), .B(N5690), .Y(N7929) );
  INVX1 gate2201 ( .A(N7903), .Y(N7930) );
  NAND2X1 gate2202 ( .A(N7903), .B(N5691), .Y(N7931) );
  NAND2X1 gate2203 ( .A(N7917), .B(N7897), .Y(N7932) );
  NAND2X1 gate2204 ( .A(N7918), .B(N7899), .Y(N7935) );
  INVX1 gate2205 ( .A(N7906), .Y(N7938) );
  NAND2X1 gate2206 ( .A(N7906), .B(N6784), .Y(N7939) );
  NAND2X1 gate2207 ( .A(N7923), .B(N7910), .Y(N7940) );
  NAND2X1 gate2208 ( .A(N6280), .B(N7924), .Y(N7943) );
  NAND2X1 gate2209 ( .A(N6292), .B(N7926), .Y(N7944) );
  NAND2X1 gate2210 ( .A(N5202), .B(N7928), .Y(N7945) );
  NAND2X1 gate2211 ( .A(N5211), .B(N7930), .Y(N7946) );
  NAND2X1 gate2212 ( .A(N6359), .B(N7938), .Y(N7951) );
  NAND2X1 gate2213 ( .A(N7943), .B(N7925), .Y(N7954) );
  NAND2X1 gate2214 ( .A(N7944), .B(N7927), .Y(N7957) );
  NAND2X1 gate2215 ( .A(N7945), .B(N7929), .Y(N7960) );
  NAND2X1 gate2216 ( .A(N7946), .B(N7931), .Y(N7963) );
  INVX1 gate2217 ( .A(N7932), .Y(N7966) );
  NAND2X1 gate2218 ( .A(N7932), .B(N6754), .Y(N7967) );
  INVX1 gate2219 ( .A(N7935), .Y(N7968) );
  NAND2X1 gate2220 ( .A(N7935), .B(N6755), .Y(N7969) );
  NAND2X1 gate2221 ( .A(N7951), .B(N7939), .Y(N7970) );
  INVX1 gate2222 ( .A(N7940), .Y(N7973) );
  NAND2X1 gate2223 ( .A(N7940), .B(N6785), .Y(N7974) );
  NAND2X1 gate2224 ( .A(N6304), .B(N7966), .Y(N7984) );
  NAND2X1 gate2225 ( .A(N6322), .B(N7968), .Y(N7985) );
  NAND2X1 gate2226 ( .A(N6370), .B(N7973), .Y(N7987) );
  AND2X1 gate2227_1 ( .A(N7957), .B(N6831), .Y(N7988_1) );
  AND2X1 gate2227 ( .A(N1157), .B(N7988_1), .Y(N7988) );
  AND2X1 gate2228_1 ( .A(N7954), .B(N6415), .Y(N7989_1) );
  AND2X1 gate2228 ( .A(N1157), .B(N7989_1), .Y(N7989) );
  AND2X1 gate2229_1 ( .A(N7957), .B(N7041), .Y(N7990_1) );
  AND2X1 gate2229 ( .A(N566), .B(N7990_1), .Y(N7990) );
  AND2X1 gate2230_1 ( .A(N7954), .B(N7177), .Y(N7991_1) );
  AND2X1 gate2230 ( .A(N566), .B(N7991_1), .Y(N7991) );
  INVX1 gate2231 ( .A(N7970), .Y(N7992) );
  NAND2X1 gate2232 ( .A(N7970), .B(N6448), .Y(N7993) );
  AND2X1 gate2233_1 ( .A(N7963), .B(N6857), .Y(N7994_1) );
  AND2X1 gate2233 ( .A(N1219), .B(N7994_1), .Y(N7994) );
  AND2X1 gate2234_1 ( .A(N7960), .B(N6441), .Y(N7995_1) );
  AND2X1 gate2234 ( .A(N1219), .B(N7995_1), .Y(N7995) );
  AND2X1 gate2235_1 ( .A(N7963), .B(N7065), .Y(N7996_1) );
  AND2X1 gate2235 ( .A(N583), .B(N7996_1), .Y(N7996) );
  AND2X1 gate2236_1 ( .A(N7960), .B(N7182), .Y(N7997_1) );
  AND2X1 gate2236 ( .A(N583), .B(N7997_1), .Y(N7997) );
  NAND2X1 gate2237 ( .A(N7984), .B(N7967), .Y(N7998) );
  NAND2X1 gate2238 ( .A(N7985), .B(N7969), .Y(N8001) );
  NAND2X1 gate2239 ( .A(N7987), .B(N7974), .Y(N8004) );
  NAND2X1 gate2240 ( .A(N6051), .B(N7992), .Y(N8009) );
  OR2X1 gate2241_1 ( .A(N7988), .B(N7989), .Y(N8013_1) );
  OR2X1 gate2241_2 ( .A(N7990), .B(N7991), .Y(N8013_2) );
  OR2X1 gate2241 ( .A(N8013_1), .B(N8013_2), .Y(N8013) );
  OR2X1 gate2242_1 ( .A(N7994), .B(N7995), .Y(N8017_1) );
  OR2X1 gate2242_2 ( .A(N7996), .B(N7997), .Y(N8017_2) );
  OR2X1 gate2242 ( .A(N8017_1), .B(N8017_2), .Y(N8017) );
  INVX1 gate2243 ( .A(N7998), .Y(N8020) );
  NAND2X1 gate2244 ( .A(N7998), .B(N6682), .Y(N8021) );
  INVX1 gate2245 ( .A(N8001), .Y(N8022) );
  NAND2X1 gate2246 ( .A(N8001), .B(N6683), .Y(N8023) );
  NAND2X1 gate2247 ( .A(N8009), .B(N7993), .Y(N8025) );
  INVX1 gate2248 ( .A(N8004), .Y(N8026) );
  NAND2X1 gate2249 ( .A(N8004), .B(N6449), .Y(N8027) );
  NAND2X1 gate2250 ( .A(N6307), .B(N8020), .Y(N8031) );
  NAND2X1 gate2251 ( .A(N6310), .B(N8022), .Y(N8032) );
  INVX1 gate2252 ( .A(N8013), .Y(N8033) );
  NAND2X1 gate2253 ( .A(N6054), .B(N8026), .Y(N8034) );
  AND2X1 gate2254 ( .A(N583), .B(N8025), .Y(N8035) );
  INVX1 gate2255 ( .A(N8017), .Y(N8036) );
  NAND2X1 gate2256 ( .A(N8031), .B(N8021), .Y(N8037) );
  NAND2X1 gate2257 ( .A(N8032), .B(N8023), .Y(N8038) );
  NAND2X1 gate2258 ( .A(N8034), .B(N8027), .Y(N8039) );
  INVX1 gate2259 ( .A(N8038), .Y(N8040) );
  AND2X1 gate2260 ( .A(N566), .B(N8037), .Y(N8041) );
  INVX1 gate2261 ( .A(N8039), .Y(N8042) );
  AND2X1 gate2262 ( .A(N8040), .B(N1157), .Y(N8043) );
  AND2X1 gate2263 ( .A(N8042), .B(N1219), .Y(N8044) );
  OR2X1 gate2264 ( .A(N8043), .B(N8041), .Y(N8045) );
  OR2X1 gate2265 ( .A(N8044), .B(N8035), .Y(N8048) );
  NAND2X1 gate2266 ( .A(N8045), .B(N8033), .Y(N8055) );
  INVX1 gate2267 ( .A(N8045), .Y(N8056) );
  NAND2X1 gate2268 ( .A(N8048), .B(N8036), .Y(N8057) );
  INVX1 gate2269 ( .A(N8048), .Y(N8058) );
  NAND2X1 gate2270 ( .A(N8013), .B(N8056), .Y(N8059) );
  NAND2X1 gate2271 ( .A(N8017), .B(N8058), .Y(N8060) );
  NAND2X1 gate2272 ( .A(N8055), .B(N8059), .Y(N8061) );
  NAND2X1 gate2273 ( .A(N8057), .B(N8060), .Y(N8064) );
  AND2X1 gate2274_1 ( .A(N8064), .B(N1777), .Y(N8071_1) );
  AND2X1 gate2274 ( .A(N3130), .B(N8071_1), .Y(N8071) );
  AND2X1 gate2275_1 ( .A(N8061), .B(N1761), .Y(N8072_1) );
  AND2X1 gate2275 ( .A(N3108), .B(N8072_1), .Y(N8072) );
  INVX1 gate2276 ( .A(N8061), .Y(N8073) );
  INVX1 gate2277 ( .A(N8064), .Y(N8074) );
  OR2X1 gate2278_1 ( .A(N7526), .B(N8071), .Y(N8075_1) );
  OR2X1 gate2278_2 ( .A(N3659), .B(N2625), .Y(N8075_2) );
  OR2X1 gate2278 ( .A(N8075_1), .B(N8075_2), .Y(N8075) );
  OR2X1 gate2279_1 ( .A(N7636), .B(N8072), .Y(N8076_1) );
  OR2X1 gate2279_2 ( .A(N3661), .B(N2627), .Y(N8076_2) );
  OR2X1 gate2279 ( .A(N8076_1), .B(N8076_2), .Y(N8076) );
  AND2X1 gate2280 ( .A(N8073), .B(N1727), .Y(N8077) );
  AND2X1 gate2281 ( .A(N8074), .B(N1727), .Y(N8078) );
  OR2X1 gate2282 ( .A(N7530), .B(N8077), .Y(N8079) );
  OR2X1 gate2283 ( .A(N7479), .B(N8078), .Y(N8082) );
  AND2X1 gate2284 ( .A(N8079), .B(N3063), .Y(N8089) );
  AND2X1 gate2285 ( .A(N8082), .B(N3063), .Y(N8090) );
  AND2X1 gate2286 ( .A(N8079), .B(N3063), .Y(N8091) );
  AND2X1 gate2287 ( .A(N8082), .B(N3063), .Y(N8092) );
  OR2X1 gate2288 ( .A(N8089), .B(N3071), .Y(N8093) );
  OR2X1 gate2289 ( .A(N8090), .B(N3072), .Y(N8096) );
  OR2X1 gate2290 ( .A(N8091), .B(N3073), .Y(N8099) );
  OR2X1 gate2291 ( .A(N8092), .B(N3074), .Y(N8102) );
  AND2X1 gate2292_1 ( .A(N8102), .B(N2779), .Y(N8113_1) );
  AND2X1 gate2292 ( .A(N2790), .B(N8113_1), .Y(N8113) );
  AND2X1 gate2293_1 ( .A(N8099), .B(N1327), .Y(N8114_1) );
  AND2X1 gate2293 ( .A(N2790), .B(N8114_1), .Y(N8114) );
  AND2X1 gate2294_1 ( .A(N8102), .B(N2801), .Y(N8115_1) );
  AND2X1 gate2294 ( .A(N2812), .B(N8115_1), .Y(N8115) );
  AND2X1 gate2295_1 ( .A(N8099), .B(N1351), .Y(N8116_1) );
  AND2X1 gate2295 ( .A(N2812), .B(N8116_1), .Y(N8116) );
  AND2X1 gate2296_1 ( .A(N8096), .B(N2681), .Y(N8117_1) );
  AND2X1 gate2296 ( .A(N2692), .B(N8117_1), .Y(N8117) );
  AND2X1 gate2297_1 ( .A(N8093), .B(N1185), .Y(N8118_1) );
  AND2X1 gate2297 ( .A(N2692), .B(N8118_1), .Y(N8118) );
  AND2X1 gate2298_1 ( .A(N8096), .B(N2756), .Y(N8119_1) );
  AND2X1 gate2298 ( .A(N2767), .B(N8119_1), .Y(N8119) );
  AND2X1 gate2299_1 ( .A(N8093), .B(N1247), .Y(N8120_1) );
  AND2X1 gate2299 ( .A(N2767), .B(N8120_1), .Y(N8120) );
  OR2X1 gate2300_1 ( .A(N8117), .B(N8118), .Y(N8121_1) );
  OR2X1 gate2300_2 ( .A(N3662), .B(N2703), .Y(N8121_2) );
  OR2X1 gate2300 ( .A(N8121_1), .B(N8121_2), .Y(N8121) );
  OR2X1 gate2301_1 ( .A(N8119), .B(N8120), .Y(N8122_1) );
  OR2X1 gate2301_2 ( .A(N3663), .B(N2778), .Y(N8122_2) );
  OR2X1 gate2301 ( .A(N8122_1), .B(N8122_2), .Y(N8122) );
  OR2X1 gate2302_1 ( .A(N8113), .B(N8114), .Y(N8123_1) );
  OR2X1 gate2302_2 ( .A(N3650), .B(N2614), .Y(N8123_2) );
  OR2X1 gate2302 ( .A(N8123_1), .B(N8123_2), .Y(N8123) );
  OR2X1 gate2303_1 ( .A(N8115), .B(N8116), .Y(N8124_1) );
  OR2X1 gate2303_2 ( .A(N3658), .B(N2622), .Y(N8124_2) );
  OR2X1 gate2303 ( .A(N8124_1), .B(N8124_2), .Y(N8124) );
  AND2X1 gate2304 ( .A(N8121), .B(N2675), .Y(N8125) );
  AND2X1 gate2305 ( .A(N8122), .B(N2750), .Y(N8126) );
  INVX1 gate2306 ( .A(N8125), .Y(N8127) );
  INVX1 gate2307 ( .A(N8126), .Y(N8128) );
endmodule



module c499_synth ( N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, 
        N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, 
        N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, 
        N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, 
        N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, 
        N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
  input N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57,
         N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109,
         N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135,
         N136, N137;
  output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734,
         N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745,
         N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
  wire   N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N293, N296, N299,
         N302, N305, N308, N311, N314, N315, N316, N317, N318, N319, N320,
         N321, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N367, N380, N393, N406,
         N419, N432, N445, N554, N555, N556, N557, N558, N559, N560, N561,
         N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572,
         N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583,
         N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594,
         N595, N596, N597, N598, N599, N600, N601, N602, N607, N620, N625,
         N630, N635, N640, N645, N650, N655, N692, N693, N694, N695, N696,
         N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N707,
         N708, N709, N710, N711, N712, N713, N714, N715, N716, N717, N718,
         N719, N720, N721, N722, N723, N594_1, N594_2, N595_1, N595_2, N596_1,
         N596_2, N597_1, N597_2, N598_1, N598_2, N599_1, N599_2, N600_1,
         N600_2, N601_1, N601_2, N602_1, N602_2, N607_1, N607_2, N620_1,
         N620_2, N620_3, N625_1, N625_2, N625_3, N630_1, N630_2, N630_3,
         N635_1, N635_2, N635_3, N640_1, N640_2, N640_3, N645_1, N645_2,
         N645_3, N650_1, N650_2, N650_3, N655_1, N655_2, N655_3;

  XOR2X1 gate1 ( .A(N1), .B(N5), .Y(N250) );
  XOR2X1 gate2 ( .A(N9), .B(N13), .Y(N251) );
  XOR2X1 gate3 ( .A(N17), .B(N21), .Y(N252) );
  XOR2X1 gate4 ( .A(N25), .B(N29), .Y(N253) );
  XOR2X1 gate5 ( .A(N33), .B(N37), .Y(N254) );
  XOR2X1 gate6 ( .A(N41), .B(N45), .Y(N255) );
  XOR2X1 gate7 ( .A(N49), .B(N53), .Y(N256) );
  XOR2X1 gate8 ( .A(N57), .B(N61), .Y(N257) );
  XOR2X1 gate9 ( .A(N65), .B(N69), .Y(N258) );
  XOR2X1 gate10 ( .A(N73), .B(N77), .Y(N259) );
  XOR2X1 gate11 ( .A(N81), .B(N85), .Y(N260) );
  XOR2X1 gate12 ( .A(N89), .B(N93), .Y(N261) );
  XOR2X1 gate13 ( .A(N97), .B(N101), .Y(N262) );
  XOR2X1 gate14 ( .A(N105), .B(N109), .Y(N263) );
  XOR2X1 gate15 ( .A(N113), .B(N117), .Y(N264) );
  XOR2X1 gate16 ( .A(N121), .B(N125), .Y(N265) );
  AND2X1 gate17 ( .A(N129), .B(N137), .Y(N266) );
  AND2X1 gate18 ( .A(N130), .B(N137), .Y(N267) );
  AND2X1 gate19 ( .A(N131), .B(N137), .Y(N268) );
  AND2X1 gate20 ( .A(N132), .B(N137), .Y(N269) );
  AND2X1 gate21 ( .A(N133), .B(N137), .Y(N270) );
  AND2X1 gate22 ( .A(N134), .B(N137), .Y(N271) );
  AND2X1 gate23 ( .A(N135), .B(N137), .Y(N272) );
  AND2X1 gate24 ( .A(N136), .B(N137), .Y(N273) );
  XOR2X1 gate25 ( .A(N1), .B(N17), .Y(N274) );
  XOR2X1 gate26 ( .A(N33), .B(N49), .Y(N275) );
  XOR2X1 gate27 ( .A(N5), .B(N21), .Y(N276) );
  XOR2X1 gate28 ( .A(N37), .B(N53), .Y(N277) );
  XOR2X1 gate29 ( .A(N9), .B(N25), .Y(N278) );
  XOR2X1 gate30 ( .A(N41), .B(N57), .Y(N279) );
  XOR2X1 gate31 ( .A(N13), .B(N29), .Y(N280) );
  XOR2X1 gate32 ( .A(N45), .B(N61), .Y(N281) );
  XOR2X1 gate33 ( .A(N65), .B(N81), .Y(N282) );
  XOR2X1 gate34 ( .A(N97), .B(N113), .Y(N283) );
  XOR2X1 gate35 ( .A(N69), .B(N85), .Y(N284) );
  XOR2X1 gate36 ( .A(N101), .B(N117), .Y(N285) );
  XOR2X1 gate37 ( .A(N73), .B(N89), .Y(N286) );
  XOR2X1 gate38 ( .A(N105), .B(N121), .Y(N287) );
  XOR2X1 gate39 ( .A(N77), .B(N93), .Y(N288) );
  XOR2X1 gate40 ( .A(N109), .B(N125), .Y(N289) );
  XOR2X1 gate41 ( .A(N250), .B(N251), .Y(N290) );
  XOR2X1 gate42 ( .A(N252), .B(N253), .Y(N293) );
  XOR2X1 gate43 ( .A(N254), .B(N255), .Y(N296) );
  XOR2X1 gate44 ( .A(N256), .B(N257), .Y(N299) );
  XOR2X1 gate45 ( .A(N258), .B(N259), .Y(N302) );
  XOR2X1 gate46 ( .A(N260), .B(N261), .Y(N305) );
  XOR2X1 gate47 ( .A(N262), .B(N263), .Y(N308) );
  XOR2X1 gate48 ( .A(N264), .B(N265), .Y(N311) );
  XOR2X1 gate49 ( .A(N274), .B(N275), .Y(N314) );
  XOR2X1 gate50 ( .A(N276), .B(N277), .Y(N315) );
  XOR2X1 gate51 ( .A(N278), .B(N279), .Y(N316) );
  XOR2X1 gate52 ( .A(N280), .B(N281), .Y(N317) );
  XOR2X1 gate53 ( .A(N282), .B(N283), .Y(N318) );
  XOR2X1 gate54 ( .A(N284), .B(N285), .Y(N319) );
  XOR2X1 gate55 ( .A(N286), .B(N287), .Y(N320) );
  XOR2X1 gate56 ( .A(N288), .B(N289), .Y(N321) );
  XOR2X1 gate57 ( .A(N290), .B(N293), .Y(N338) );
  XOR2X1 gate58 ( .A(N296), .B(N299), .Y(N339) );
  XOR2X1 gate59 ( .A(N290), .B(N296), .Y(N340) );
  XOR2X1 gate60 ( .A(N293), .B(N299), .Y(N341) );
  XOR2X1 gate61 ( .A(N302), .B(N305), .Y(N342) );
  XOR2X1 gate62 ( .A(N308), .B(N311), .Y(N343) );
  XOR2X1 gate63 ( .A(N302), .B(N308), .Y(N344) );
  XOR2X1 gate64 ( .A(N305), .B(N311), .Y(N345) );
  XOR2X1 gate65 ( .A(N266), .B(N342), .Y(N346) );
  XOR2X1 gate66 ( .A(N267), .B(N343), .Y(N347) );
  XOR2X1 gate67 ( .A(N268), .B(N344), .Y(N348) );
  XOR2X1 gate68 ( .A(N269), .B(N345), .Y(N349) );
  XOR2X1 gate69 ( .A(N270), .B(N338), .Y(N350) );
  XOR2X1 gate70 ( .A(N271), .B(N339), .Y(N351) );
  XOR2X1 gate71 ( .A(N272), .B(N340), .Y(N352) );
  XOR2X1 gate72 ( .A(N273), .B(N341), .Y(N353) );
  XOR2X1 gate73 ( .A(N314), .B(N346), .Y(N354) );
  XOR2X1 gate74 ( .A(N315), .B(N347), .Y(N367) );
  XOR2X1 gate75 ( .A(N316), .B(N348), .Y(N380) );
  XOR2X1 gate76 ( .A(N317), .B(N349), .Y(N393) );
  XOR2X1 gate77 ( .A(N318), .B(N350), .Y(N406) );
  XOR2X1 gate78 ( .A(N319), .B(N351), .Y(N419) );
  XOR2X1 gate79 ( .A(N320), .B(N352), .Y(N432) );
  XOR2X1 gate80 ( .A(N321), .B(N353), .Y(N445) );
  INVX1 gate81 ( .A(N354), .Y(N554) );
  INVX1 gate82 ( .A(N367), .Y(N555) );
  INVX1 gate83 ( .A(N380), .Y(N556) );
  INVX1 gate84 ( .A(N354), .Y(N557) );
  INVX1 gate85 ( .A(N367), .Y(N558) );
  INVX1 gate86 ( .A(N393), .Y(N559) );
  INVX1 gate87 ( .A(N354), .Y(N560) );
  INVX1 gate88 ( .A(N380), .Y(N561) );
  INVX1 gate89 ( .A(N393), .Y(N562) );
  INVX1 gate90 ( .A(N367), .Y(N563) );
  INVX1 gate91 ( .A(N380), .Y(N564) );
  INVX1 gate92 ( .A(N393), .Y(N565) );
  INVX1 gate93 ( .A(N419), .Y(N566) );
  INVX1 gate94 ( .A(N445), .Y(N567) );
  INVX1 gate95 ( .A(N419), .Y(N568) );
  INVX1 gate96 ( .A(N432), .Y(N569) );
  INVX1 gate97 ( .A(N406), .Y(N570) );
  INVX1 gate98 ( .A(N445), .Y(N571) );
  INVX1 gate99 ( .A(N406), .Y(N572) );
  INVX1 gate100 ( .A(N432), .Y(N573) );
  INVX1 gate101 ( .A(N406), .Y(N574) );
  INVX1 gate102 ( .A(N419), .Y(N575) );
  INVX1 gate103 ( .A(N432), .Y(N576) );
  INVX1 gate104 ( .A(N406), .Y(N577) );
  INVX1 gate105 ( .A(N419), .Y(N578) );
  INVX1 gate106 ( .A(N445), .Y(N579) );
  INVX1 gate107 ( .A(N406), .Y(N580) );
  INVX1 gate108 ( .A(N432), .Y(N581) );
  INVX1 gate109 ( .A(N445), .Y(N582) );
  INVX1 gate110 ( .A(N419), .Y(N583) );
  INVX1 gate111 ( .A(N432), .Y(N584) );
  INVX1 gate112 ( .A(N445), .Y(N585) );
  INVX1 gate113 ( .A(N367), .Y(N586) );
  INVX1 gate114 ( .A(N393), .Y(N587) );
  INVX1 gate115 ( .A(N367), .Y(N588) );
  INVX1 gate116 ( .A(N380), .Y(N589) );
  INVX1 gate117 ( .A(N354), .Y(N590) );
  INVX1 gate118 ( .A(N393), .Y(N591) );
  INVX1 gate119 ( .A(N354), .Y(N592) );
  INVX1 gate120 ( .A(N380), .Y(N593) );
  AND2X1 gate121_1 ( .A(N554), .B(N555), .Y(N594_1) );
  AND2X1 gate121_2 ( .A(N556), .B(N393), .Y(N594_2) );
  AND2X1 gate121 ( .A(N594_1), .B(N594_2), .Y(N594) );
  AND2X1 gate122_1 ( .A(N557), .B(N558), .Y(N595_1) );
  AND2X1 gate122_2 ( .A(N380), .B(N559), .Y(N595_2) );
  AND2X1 gate122 ( .A(N595_1), .B(N595_2), .Y(N595) );
  AND2X1 gate123_1 ( .A(N560), .B(N367), .Y(N596_1) );
  AND2X1 gate123_2 ( .A(N561), .B(N562), .Y(N596_2) );
  AND2X1 gate123 ( .A(N596_1), .B(N596_2), .Y(N596) );
  AND2X1 gate124_1 ( .A(N354), .B(N563), .Y(N597_1) );
  AND2X1 gate124_2 ( .A(N564), .B(N565), .Y(N597_2) );
  AND2X1 gate124 ( .A(N597_1), .B(N597_2), .Y(N597) );
  AND2X1 gate125_1 ( .A(N574), .B(N575), .Y(N598_1) );
  AND2X1 gate125_2 ( .A(N576), .B(N445), .Y(N598_2) );
  AND2X1 gate125 ( .A(N598_1), .B(N598_2), .Y(N598) );
  AND2X1 gate126_1 ( .A(N577), .B(N578), .Y(N599_1) );
  AND2X1 gate126_2 ( .A(N432), .B(N579), .Y(N599_2) );
  AND2X1 gate126 ( .A(N599_1), .B(N599_2), .Y(N599) );
  AND2X1 gate127_1 ( .A(N580), .B(N419), .Y(N600_1) );
  AND2X1 gate127_2 ( .A(N581), .B(N582), .Y(N600_2) );
  AND2X1 gate127 ( .A(N600_1), .B(N600_2), .Y(N600) );
  AND2X1 gate128_1 ( .A(N406), .B(N583), .Y(N601_1) );
  AND2X1 gate128_2 ( .A(N584), .B(N585), .Y(N601_2) );
  AND2X1 gate128 ( .A(N601_1), .B(N601_2), .Y(N601) );
  OR2X1 gate129_1 ( .A(N594), .B(N595), .Y(N602_1) );
  OR2X1 gate129_2 ( .A(N596), .B(N597), .Y(N602_2) );
  OR2X1 gate129 ( .A(N602_1), .B(N602_2), .Y(N602) );
  OR2X1 gate130_1 ( .A(N598), .B(N599), .Y(N607_1) );
  OR2X1 gate130_2 ( .A(N600), .B(N601), .Y(N607_2) );
  OR2X1 gate130 ( .A(N607_1), .B(N607_2), .Y(N607) );
  AND2X1 gate131_1 ( .A(N406), .B(N566), .Y(N620_1) );
  AND2X1 gate131_2 ( .A(N432), .B(N567), .Y(N620_2) );
  AND2X1 gate131_3 ( .A(N602), .B(N620_1), .Y(N620_3) );
  AND2X1 gate131 ( .A(N620_2), .B(N620_3), .Y(N620) );
  AND2X1 gate132_1 ( .A(N406), .B(N568), .Y(N625_1) );
  AND2X1 gate132_2 ( .A(N569), .B(N445), .Y(N625_2) );
  AND2X1 gate132_3 ( .A(N602), .B(N625_1), .Y(N625_3) );
  AND2X1 gate132 ( .A(N625_2), .B(N625_3), .Y(N625) );
  AND2X1 gate133_1 ( .A(N570), .B(N419), .Y(N630_1) );
  AND2X1 gate133_2 ( .A(N432), .B(N571), .Y(N630_2) );
  AND2X1 gate133_3 ( .A(N602), .B(N630_1), .Y(N630_3) );
  AND2X1 gate133 ( .A(N630_2), .B(N630_3), .Y(N630) );
  AND2X1 gate134_1 ( .A(N572), .B(N419), .Y(N635_1) );
  AND2X1 gate134_2 ( .A(N573), .B(N445), .Y(N635_2) );
  AND2X1 gate134_3 ( .A(N602), .B(N635_1), .Y(N635_3) );
  AND2X1 gate134 ( .A(N635_2), .B(N635_3), .Y(N635) );
  AND2X1 gate135_1 ( .A(N354), .B(N586), .Y(N640_1) );
  AND2X1 gate135_2 ( .A(N380), .B(N587), .Y(N640_2) );
  AND2X1 gate135_3 ( .A(N607), .B(N640_1), .Y(N640_3) );
  AND2X1 gate135 ( .A(N640_2), .B(N640_3), .Y(N640) );
  AND2X1 gate136_1 ( .A(N354), .B(N588), .Y(N645_1) );
  AND2X1 gate136_2 ( .A(N589), .B(N393), .Y(N645_2) );
  AND2X1 gate136_3 ( .A(N607), .B(N645_1), .Y(N645_3) );
  AND2X1 gate136 ( .A(N645_2), .B(N645_3), .Y(N645) );
  AND2X1 gate137_1 ( .A(N590), .B(N367), .Y(N650_1) );
  AND2X1 gate137_2 ( .A(N380), .B(N591), .Y(N650_2) );
  AND2X1 gate137_3 ( .A(N607), .B(N650_1), .Y(N650_3) );
  AND2X1 gate137 ( .A(N650_2), .B(N650_3), .Y(N650) );
  AND2X1 gate138_1 ( .A(N592), .B(N367), .Y(N655_1) );
  AND2X1 gate138_2 ( .A(N593), .B(N393), .Y(N655_2) );
  AND2X1 gate138_3 ( .A(N607), .B(N655_1), .Y(N655_3) );
  AND2X1 gate138 ( .A(N655_2), .B(N655_3), .Y(N655) );
  AND2X1 gate139 ( .A(N354), .B(N620), .Y(N692) );
  AND2X1 gate140 ( .A(N367), .B(N620), .Y(N693) );
  AND2X1 gate141 ( .A(N380), .B(N620), .Y(N694) );
  AND2X1 gate142 ( .A(N393), .B(N620), .Y(N695) );
  AND2X1 gate143 ( .A(N354), .B(N625), .Y(N696) );
  AND2X1 gate144 ( .A(N367), .B(N625), .Y(N697) );
  AND2X1 gate145 ( .A(N380), .B(N625), .Y(N698) );
  AND2X1 gate146 ( .A(N393), .B(N625), .Y(N699) );
  AND2X1 gate147 ( .A(N354), .B(N630), .Y(N700) );
  AND2X1 gate148 ( .A(N367), .B(N630), .Y(N701) );
  AND2X1 gate149 ( .A(N380), .B(N630), .Y(N702) );
  AND2X1 gate150 ( .A(N393), .B(N630), .Y(N703) );
  AND2X1 gate151 ( .A(N354), .B(N635), .Y(N704) );
  AND2X1 gate152 ( .A(N367), .B(N635), .Y(N705) );
  AND2X1 gate153 ( .A(N380), .B(N635), .Y(N706) );
  AND2X1 gate154 ( .A(N393), .B(N635), .Y(N707) );
  AND2X1 gate155 ( .A(N406), .B(N640), .Y(N708) );
  AND2X1 gate156 ( .A(N419), .B(N640), .Y(N709) );
  AND2X1 gate157 ( .A(N432), .B(N640), .Y(N710) );
  AND2X1 gate158 ( .A(N445), .B(N640), .Y(N711) );
  AND2X1 gate159 ( .A(N406), .B(N645), .Y(N712) );
  AND2X1 gate160 ( .A(N419), .B(N645), .Y(N713) );
  AND2X1 gate161 ( .A(N432), .B(N645), .Y(N714) );
  AND2X1 gate162 ( .A(N445), .B(N645), .Y(N715) );
  AND2X1 gate163 ( .A(N406), .B(N650), .Y(N716) );
  AND2X1 gate164 ( .A(N419), .B(N650), .Y(N717) );
  AND2X1 gate165 ( .A(N432), .B(N650), .Y(N718) );
  AND2X1 gate166 ( .A(N445), .B(N650), .Y(N719) );
  AND2X1 gate167 ( .A(N406), .B(N655), .Y(N720) );
  AND2X1 gate168 ( .A(N419), .B(N655), .Y(N721) );
  AND2X1 gate169 ( .A(N432), .B(N655), .Y(N722) );
  AND2X1 gate170 ( .A(N445), .B(N655), .Y(N723) );
  XOR2X1 gate171 ( .A(N1), .B(N692), .Y(N724) );
  XOR2X1 gate172 ( .A(N5), .B(N693), .Y(N725) );
  XOR2X1 gate173 ( .A(N9), .B(N694), .Y(N726) );
  XOR2X1 gate174 ( .A(N13), .B(N695), .Y(N727) );
  XOR2X1 gate175 ( .A(N17), .B(N696), .Y(N728) );
  XOR2X1 gate176 ( .A(N21), .B(N697), .Y(N729) );
  XOR2X1 gate177 ( .A(N25), .B(N698), .Y(N730) );
  XOR2X1 gate178 ( .A(N29), .B(N699), .Y(N731) );
  XOR2X1 gate179 ( .A(N33), .B(N700), .Y(N732) );
  XOR2X1 gate180 ( .A(N37), .B(N701), .Y(N733) );
  XOR2X1 gate181 ( .A(N41), .B(N702), .Y(N734) );
  XOR2X1 gate182 ( .A(N45), .B(N703), .Y(N735) );
  XOR2X1 gate183 ( .A(N49), .B(N704), .Y(N736) );
  XOR2X1 gate184 ( .A(N53), .B(N705), .Y(N737) );
  XOR2X1 gate185 ( .A(N57), .B(N706), .Y(N738) );
  XOR2X1 gate186 ( .A(N61), .B(N707), .Y(N739) );
  XOR2X1 gate187 ( .A(N65), .B(N708), .Y(N740) );
  XOR2X1 gate188 ( .A(N69), .B(N709), .Y(N741) );
  XOR2X1 gate189 ( .A(N73), .B(N710), .Y(N742) );
  XOR2X1 gate190 ( .A(N77), .B(N711), .Y(N743) );
  XOR2X1 gate191 ( .A(N81), .B(N712), .Y(N744) );
  XOR2X1 gate192 ( .A(N85), .B(N713), .Y(N745) );
  XOR2X1 gate193 ( .A(N89), .B(N714), .Y(N746) );
  XOR2X1 gate194 ( .A(N93), .B(N715), .Y(N747) );
  XOR2X1 gate195 ( .A(N97), .B(N716), .Y(N748) );
  XOR2X1 gate196 ( .A(N101), .B(N717), .Y(N749) );
  XOR2X1 gate197 ( .A(N105), .B(N718), .Y(N750) );
  XOR2X1 gate198 ( .A(N109), .B(N719), .Y(N751) );
  XOR2X1 gate199 ( .A(N113), .B(N720), .Y(N752) );
  XOR2X1 gate200 ( .A(N117), .B(N721), .Y(N753) );
  XOR2X1 gate201 ( .A(N121), .B(N722), .Y(N754) );
  XOR2X1 gate202 ( .A(N125), .B(N723), .Y(N755) );
endmodule


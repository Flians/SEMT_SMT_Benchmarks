
module c7552_synth ( N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, 
        N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, 
        N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, 
        N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, 
        N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, 
        N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, 
        N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, 
        N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, 
        N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, 
        N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, 
        N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, 
        N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, 
        N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, 
        N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, 
        N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, 
        N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, 
        N346, N349, N352, N355, N358, N361, N364, N367, N382, N241_I, N387, 
        N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, 
        N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, 
        N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, 
        N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, 
        N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, 
        N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, 
        N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, 
        N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, 
        N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, 
        N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, 
        N10908, N11333, N11334, N11340, N11342, N241_O );
  input N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47,
         N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110,
         N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133,
         N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245,
         N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280,
         N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316,
         N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349,
         N352, N355, N358, N361, N364, N367, N382, N241_I;
  output N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507,
         N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543,
         N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567,
         N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884,
         N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490,
         N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111,
         N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576,
         N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713,
         N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760,
         N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840,
         N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908,
         N11333, N11334, N11340, N11342, N241_O;
  wire   N467, N469, N494, N528, N575, N578, N585, N590, N593, N596, N599,
         N604, N609, N614, N625, N628, N632, N636, N641, N642, N644, N651,
         N657, N660, N666, N672, N673, N674, N676, N682, N688, N689, N695,
         N700, N705, N706, N708, N715, N721, N727, N733, N734, N742, N748,
         N749, N750, N758, N759, N762, N768, N774, N780, N786, N794, N800,
         N806, N812, N814, N821, N827, N833, N839, N845, N853, N859, N865,
         N871, N886, N887, N957, N1028, N1029, N1109, N1115, N1116, N1119,
         N1125, N1132, N1136, N1141, N1147, N1154, N1160, N1167, N1174, N1175,
         N1182, N1189, N1194, N1199, N1206, N1211, N1218, N1222, N1227, N1233,
         N1240, N1244, N1249, N1256, N1263, N1270, N1277, N1284, N1287, N1290,
         N1293, N1296, N1299, N1302, N1305, N1308, N1311, N1314, N1317, N1320,
         N1323, N1326, N1329, N1332, N1335, N1338, N1341, N1344, N1347, N1350,
         N1353, N1356, N1359, N1362, N1365, N1368, N1371, N1374, N1377, N1380,
         N1383, N1386, N1389, N1392, N1395, N1398, N1401, N1404, N1407, N1410,
         N1413, N1416, N1419, N1422, N1425, N1428, N1431, N1434, N1437, N1440,
         N1443, N1446, N1449, N1452, N1455, N1458, N1461, N1464, N1467, N1470,
         N1473, N1476, N1479, N1482, N1485, N1537, N1551, N1649, N1703, N1708,
         N1713, N1721, N1758, N1782, N1783, N1789, N1793, N1794, N1795, N1796,
         N1797, N1798, N1799, N1805, N1811, N1812, N1813, N1814, N1815, N1816,
         N1817, N1818, N1819, N1820, N1821, N1822, N1828, N1829, N1830, N1832,
         N1833, N1834, N1835, N1839, N1840, N1841, N1842, N1843, N1845, N1851,
         N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864, N1865, N1866,
         N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874, N1875, N1876,
         N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884, N1885, N1892,
         N1899, N1906, N1913, N1919, N1926, N1927, N1928, N1929, N1930, N1931,
         N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941,
         N1942, N1943, N1944, N1945, N1946, N1947, N1953, N1957, N1958, N1959,
         N1960, N1961, N1962, N1963, N1965, N1966, N1967, N1968, N1969, N1970,
         N1971, N1972, N1973, N1974, N1975, N1976, N1977, N1983, N1989, N1990,
         N1991, N1992, N1993, N1994, N1995, N1996, N1997, N2003, N2010, N2011,
         N2012, N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021,
         N2022, N2023, N2024, N2031, N2038, N2045, N2052, N2058, N2064, N2065,
         N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073, N2074, N2081,
         N2086, N2107, N2108, N2110, N2111, N2112, N2113, N2114, N2115, N2117,
         N2171, N2172, N2230, N2231, N2235, N2239, N2240, N2241, N2242, N2243,
         N2244, N2245, N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253,
         N2254, N2255, N2256, N2257, N2267, N2268, N2269, N2274, N2275, N2277,
         N2278, N2279, N2280, N2281, N2282, N2283, N2284, N2285, N2286, N2287,
         N2293, N2299, N2300, N2301, N2302, N2303, N2304, N2305, N2306, N2307,
         N2308, N2309, N2315, N2321, N2322, N2323, N2324, N2325, N2326, N2327,
         N2328, N2329, N2330, N2331, N2337, N2338, N2339, N2340, N2341, N2342,
         N2343, N2344, N2345, N2346, N2347, N2348, N2349, N2350, N2351, N2352,
         N2353, N2354, N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362,
         N2363, N2364, N2365, N2366, N2367, N2368, N2374, N2375, N2376, N2377,
         N2378, N2379, N2380, N2381, N2382, N2383, N2384, N2390, N2396, N2397,
         N2398, N2399, N2400, N2401, N2402, N2403, N2404, N2405, N2406, N2412,
         N2418, N2419, N2420, N2421, N2422, N2423, N2424, N2425, N2426, N2427,
         N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2435, N2436, N2437,
         N2441, N2442, N2446, N2450, N2454, N2458, N2462, N2466, N2470, N2474,
         N2478, N2482, N2488, N2496, N2502, N2508, N2523, N2533, N2537, N2538,
         N2542, N2546, N2550, N2554, N2561, N2567, N2573, N2604, N2607, N2611,
         N2615, N2619, N2626, N2632, N2638, N2644, N2650, N2653, N2654, N2658,
         N2662, N2666, N2670, N2674, N2680, N2688, N2692, N2696, N2700, N2704,
         N2728, N2729, N2733, N2737, N2741, N2745, N2749, N2753, N2757, N2761,
         N2765, N2766, N2769, N2772, N2775, N2778, N2781, N2784, N2787, N2790,
         N2793, N2796, N2866, N2867, N2868, N2869, N2878, N2913, N2914, N2915,
         N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925,
         N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935,
         N2936, N2937, N2988, N3005, N3006, N3007, N3008, N3009, N3020, N3021,
         N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3032, N3033,
         N3034, N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3061, N3064,
         N3067, N3070, N3073, N3080, N3096, N3097, N3101, N3107, N3114, N3122,
         N3126, N3130, N3131, N3134, N3135, N3136, N3137, N3140, N3144, N3149,
         N3155, N3159, N3167, N3168, N3169, N3173, N3178, N3184, N3185, N3189,
         N3195, N3202, N3210, N3211, N3215, N3221, N3228, N3229, N3232, N3236,
         N3241, N3247, N3251, N3255, N3259, N3263, N3267, N3273, N3281, N3287,
         N3293, N3299, N3303, N3307, N3311, N3315, N3322, N3328, N3334, N3340,
         N3343, N3349, N3355, N3361, N3362, N3363, N3364, N3365, N3366, N3367,
         N3368, N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3379, N3380,
         N3381, N3384, N3390, N3398, N3404, N3410, N3416, N3420, N3424, N3428,
         N3432, N3436, N3440, N3444, N3448, N3452, N3453, N3454, N3458, N3462,
         N3466, N3470, N3474, N3478, N3482, N3486, N3487, N3490, N3493, N3496,
         N3499, N3502, N3507, N3510, N3515, N3518, N3521, N3524, N3527, N3530,
         N3535, N3539, N3542, N3545, N3548, N3551, N3552, N3553, N3557, N3560,
         N3563, N3566, N3569, N3570, N3571, N3574, N3577, N3580, N3583, N3586,
         N3589, N3592, N3595, N3598, N3601, N3604, N3607, N3610, N3613, N3616,
         N3619, N3622, N3625, N3628, N3631, N3634, N3637, N3640, N3643, N3646,
         N3649, N3652, N3655, N3658, N3661, N3664, N3667, N3670, N3673, N3676,
         N3679, N3682, N3685, N3688, N3691, N3694, N3697, N3700, N3703, N3706,
         N3709, N3712, N3715, N3718, N3721, N3724, N3727, N3730, N3733, N3736,
         N3739, N3742, N3745, N3748, N3751, N3754, N3757, N3760, N3763, N3766,
         N3769, N3772, N3775, N3778, N3781, N3782, N3783, N3786, N3789, N3792,
         N3795, N3798, N3801, N3804, N3807, N3810, N3813, N3816, N3819, N3822,
         N3825, N3828, N3831, N3834, N3837, N3840, N3843, N3846, N3849, N3852,
         N3855, N3858, N3861, N3864, N3867, N3870, N3873, N3876, N3879, N3882,
         N3885, N3888, N3891, N3953, N3954, N3955, N3956, N3958, N3964, N4193,
         N4303, N4308, N4313, N4326, N4327, N4333, N4334, N4411, N4412, N4463,
         N4464, N4465, N4466, N4467, N4468, N4469, N4470, N4471, N4472, N4473,
         N4474, N4475, N4476, N4477, N4478, N4479, N4480, N4481, N4482, N4483,
         N4484, N4485, N4486, N4487, N4488, N4489, N4490, N4491, N4492, N4493,
         N4494, N4495, N4496, N4497, N4498, N4499, N4500, N4501, N4502, N4503,
         N4504, N4505, N4506, N4507, N4508, N4509, N4510, N4511, N4512, N4513,
         N4514, N4515, N4516, N4517, N4518, N4519, N4520, N4521, N4522, N4523,
         N4524, N4525, N4526, N4527, N4528, N4529, N4530, N4531, N4532, N4533,
         N4534, N4535, N4536, N4537, N4538, N4539, N4540, N4541, N4542, N4543,
         N4544, N4545, N4549, N4555, N4562, N4563, N4566, N4570, N4575, N4576,
         N4577, N4581, N4586, N4592, N4593, N4597, N4603, N4610, N4611, N4612,
         N4613, N4614, N4615, N4616, N4617, N4618, N4619, N4620, N4621, N4622,
         N4623, N4624, N4625, N4626, N4627, N4628, N4629, N4630, N4631, N4632,
         N4633, N4634, N4635, N4636, N4637, N4638, N4639, N4640, N4641, N4642,
         N4643, N4644, N4645, N4646, N4647, N4648, N4649, N4650, N4651, N4652,
         N4653, N4656, N4657, N4661, N4667, N4674, N4675, N4678, N4682, N4687,
         N4693, N4694, N4695, N4696, N4697, N4698, N4699, N4700, N4701, N4702,
         N4706, N4711, N4717, N4718, N4722, N4728, N4735, N4743, N4744, N4745,
         N4746, N4747, N4748, N4749, N4750, N4751, N4752, N4753, N4754, N4755,
         N4756, N4757, N4758, N4759, N4760, N4761, N4762, N4763, N4764, N4765,
         N4766, N4767, N4768, N4769, N4775, N4776, N4777, N4778, N4779, N4780,
         N4781, N4782, N4783, N4784, N4789, N4790, N4793, N4794, N4795, N4796,
         N4799, N4800, N4801, N4802, N4803, N4806, N4809, N4810, N4813, N4814,
         N4817, N4820, N4823, N4826, N4829, N4832, N4835, N4838, N4841, N4844,
         N4847, N4850, N4853, N4856, N4859, N4862, N4865, N4868, N4871, N4874,
         N4877, N4880, N4883, N4886, N4889, N4892, N4895, N4898, N4901, N4904,
         N4907, N4910, N4913, N4916, N4919, N4922, N4925, N4928, N4931, N4934,
         N4937, N4940, N4943, N4946, N4949, N4952, N4955, N4958, N4961, N4964,
         N4967, N4970, N4973, N4976, N4979, N4982, N4985, N4988, N4991, N4994,
         N4997, N5000, N5003, N5006, N5009, N5012, N5015, N5018, N5021, N5024,
         N5027, N5030, N5033, N5036, N5039, N5042, N5045, N5046, N5047, N5048,
         N5049, N5052, N5055, N5058, N5061, N5064, N5065, N5066, N5067, N5068,
         N5071, N5074, N5077, N5080, N5083, N5086, N5089, N5092, N5095, N5098,
         N5101, N5104, N5107, N5110, N5111, N5112, N5113, N5114, N5117, N5120,
         N5123, N5126, N5129, N5132, N5135, N5138, N5141, N5144, N5147, N5150,
         N5153, N5156, N5159, N5162, N5165, N5166, N5167, N5168, N5169, N5170,
         N5171, N5172, N5173, N5174, N5175, N5176, N5177, N5178, N5179, N5180,
         N5181, N5182, N5183, N5184, N5185, N5186, N5187, N5188, N5189, N5190,
         N5191, N5192, N5193, N5196, N5197, N5198, N5199, N5200, N5201, N5202,
         N5203, N5204, N5205, N5206, N5207, N5208, N5209, N5210, N5211, N5212,
         N5213, N5283, N5284, N5285, N5286, N5287, N5288, N5289, N5290, N5291,
         N5292, N5293, N5294, N5295, N5296, N5297, N5298, N5299, N5300, N5314,
         N5315, N5316, N5317, N5318, N5319, N5320, N5321, N5322, N5323, N5324,
         N5363, N5364, N5365, N5366, N5367, N5425, N5426, N5427, N5429, N5430,
         N5431, N5432, N5433, N5451, N5452, N5453, N5454, N5455, N5456, N5457,
         N5469, N5474, N5475, N5476, N5477, N5571, N5572, N5573, N5574, N5584,
         N5585, N5586, N5587, N5602, N5603, N5604, N5605, N5631, N5632, N5640,
         N5654, N5670, N5683, N5690, N5697, N5707, N5718, N5728, N5735, N5736,
         N5740, N5744, N5747, N5751, N5755, N5758, N5762, N5766, N5769, N5770,
         N5771, N5778, N5789, N5799, N5807, N5821, N5837, N5850, N5856, N5863,
         N5870, N5881, N5892, N5898, N5905, N5915, N5926, N5936, N5943, N5944,
         N5945, N5946, N5947, N5948, N5949, N5950, N5951, N5952, N5953, N5954,
         N5955, N5956, N5957, N5958, N5959, N5960, N5966, N5967, N5968, N5969,
         N5970, N5971, N5972, N5973, N5974, N5975, N5976, N5977, N5978, N5979,
         N5980, N5981, N5989, N5990, N5991, N5996, N6000, N6003, N6009, N6014,
         N6018, N6021, N6022, N6023, N6024, N6025, N6026, N6027, N6028, N6029,
         N6030, N6031, N6032, N6033, N6034, N6035, N6036, N6037, N6038, N6039,
         N6040, N6041, N6047, N6052, N6056, N6059, N6060, N6061, N6062, N6063,
         N6064, N6065, N6066, N6067, N6068, N6069, N6070, N6071, N6072, N6073,
         N6074, N6075, N6076, N6077, N6078, N6079, N6083, N6087, N6090, N6091,
         N6092, N6093, N6094, N6095, N6096, N6097, N6098, N6099, N6100, N6101,
         N6102, N6103, N6104, N6105, N6106, N6107, N6108, N6109, N6110, N6111,
         N6112, N6113, N6114, N6115, N6116, N6117, N6118, N6119, N6120, N6121,
         N6122, N6123, N6124, N6125, N6126, N6127, N6131, N6135, N6136, N6137,
         N6141, N6145, N6148, N6149, N6150, N6151, N6152, N6153, N6154, N6155,
         N6156, N6157, N6158, N6159, N6160, N6161, N6162, N6163, N6164, N6165,
         N6166, N6170, N6174, N6177, N6181, N6182, N6183, N6184, N6185, N6186,
         N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6195, N6196,
         N6199, N6202, N6203, N6204, N6207, N6210, N6213, N6214, N6217, N6220,
         N6223, N6224, N6225, N6226, N6227, N6228, N6229, N6230, N6231, N6232,
         N6235, N6236, N6239, N6240, N6241, N6242, N6243, N6246, N6249, N6252,
         N6255, N6256, N6257, N6258, N6259, N6260, N6261, N6262, N6263, N6266,
         N6540, N6541, N6542, N6543, N6544, N6545, N6546, N6547, N6555, N6556,
         N6557, N6558, N6559, N6560, N6561, N6569, N6594, N6595, N6596, N6597,
         N6598, N6599, N6600, N6601, N6602, N6603, N6604, N6605, N6606, N6621,
         N6622, N6623, N6624, N6625, N6626, N6627, N6628, N6629, N6639, N6640,
         N6641, N6642, N6643, N6644, N6645, N6646, N6647, N6648, N6649, N6650,
         N6651, N6652, N6653, N6654, N6655, N6656, N6657, N6658, N6659, N6660,
         N6661, N6668, N6677, N6678, N6679, N6680, N6681, N6682, N6683, N6684,
         N6685, N6686, N6687, N6688, N6689, N6690, N6702, N6703, N6704, N6705,
         N6706, N6707, N6708, N6709, N6710, N6711, N6712, N6729, N6730, N6731,
         N6732, N6733, N6734, N6735, N6736, N6741, N6742, N6743, N6744, N6751,
         N6752, N6753, N6754, N6755, N6756, N6757, N6758, N6761, N6762, N6766,
         N6767, N6768, N6769, N6770, N6771, N6772, N6773, N6774, N6775, N6776,
         N6777, N6778, N6779, N6780, N6781, N6782, N6783, N6784, N6787, N6788,
         N6789, N6790, N6791, N6792, N6793, N6794, N6795, N6796, N6797, N6800,
         N6803, N6806, N6809, N6812, N6815, N6818, N6821, N6824, N6827, N6830,
         N6833, N6836, N6837, N6838, N6839, N6840, N6841, N6842, N6843, N6844,
         N6845, N6848, N6849, N6850, N6851, N6852, N6853, N6854, N6855, N6856,
         N6857, N6858, N6859, N6860, N6861, N6862, N6863, N6864, N6865, N6866,
         N6867, N6870, N6871, N6872, N6873, N6874, N6875, N6876, N6877, N6878,
         N6879, N6880, N6881, N6884, N6885, N6886, N6887, N6888, N6889, N6890,
         N6891, N6892, N6893, N6894, N6901, N6912, N6923, N6929, N6936, N6946,
         N6957, N6967, N6968, N6969, N6970, N6977, N6988, N6998, N7006, N7020,
         N7036, N7049, N7055, N7056, N7057, N7060, N7061, N7062, N7063, N7064,
         N7065, N7066, N7067, N7068, N7073, N7077, N7080, N7086, N7091, N7095,
         N7098, N7099, N7100, N7103, N7104, N7105, N7106, N7107, N7114, N7125,
         N7136, N7142, N7149, N7159, N7170, N7180, N7187, N7188, N7191, N7194,
         N7198, N7202, N7205, N7209, N7213, N7216, N7219, N7222, N7229, N7240,
         N7250, N7258, N7272, N7288, N7301, N7307, N7314, N7318, N7322, N7325,
         N7328, N7331, N7334, N7337, N7340, N7343, N7346, N7351, N7355, N7358,
         N7364, N7369, N7373, N7376, N7377, N7378, N7381, N7384, N7387, N7391,
         N7394, N7398, N7402, N7405, N7408, N7411, N7414, N7417, N7420, N7423,
         N7426, N7429, N7432, N7435, N7438, N7441, N7444, N7447, N7450, N7453,
         N7456, N7459, N7462, N7465, N7468, N7471, N7474, N7477, N7478, N7479,
         N7482, N7485, N7488, N7491, N7494, N7497, N7500, N7503, N7506, N7509,
         N7512, N7515, N7518, N7521, N7524, N7527, N7530, N7533, N7536, N7539,
         N7542, N7545, N7548, N7551, N7552, N7553, N7556, N7557, N7558, N7559,
         N7560, N7563, N7566, N7569, N7572, N7573, N7574, N7577, N7580, N7581,
         N7582, N7585, N7588, N7591, N7609, N7613, N7620, N7649, N7650, N7655,
         N7659, N7668, N7671, N7744, N7822, N7825, N7826, N7852, N8114, N8117,
         N8131, N8134, N8144, N8145, N8146, N8156, N8166, N8169, N8183, N8186,
         N8196, N8200, N8204, N8208, N8216, N8217, N8218, N8219, N8232, N8233,
         N8242, N8243, N8244, N8245, N8246, N8247, N8248, N8249, N8250, N8251,
         N8252, N8253, N8254, N8260, N8261, N8262, N8269, N8274, N8275, N8276,
         N8277, N8278, N8279, N8280, N8281, N8282, N8283, N8284, N8285, N8288,
         N8294, N8295, N8296, N8297, N8298, N8307, N8315, N8317, N8319, N8321,
         N8322, N8323, N8324, N8325, N8326, N8333, N8337, N8338, N8339, N8340,
         N8341, N8342, N8343, N8344, N8345, N8346, N8347, N8348, N8349, N8350,
         N8351, N8352, N8353, N8354, N8355, N8356, N8357, N8358, N8365, N8369,
         N8370, N8371, N8372, N8373, N8374, N8375, N8376, N8377, N8378, N8379,
         N8380, N8381, N8382, N8383, N8384, N8385, N8386, N8387, N8388, N8389,
         N8390, N8391, N8392, N8393, N8394, N8404, N8405, N8409, N8410, N8411,
         N8412, N8415, N8416, N8417, N8418, N8421, N8430, N8433, N8434, N8435,
         N8436, N8437, N8438, N8439, N8440, N8441, N8442, N8443, N8444, N8447,
         N8448, N8449, N8450, N8451, N8452, N8453, N8454, N8455, N8456, N8457,
         N8460, N8463, N8466, N8469, N8470, N8471, N8474, N8477, N8480, N8483,
         N8484, N8485, N8488, N8489, N8490, N8491, N8492, N8493, N8494, N8495,
         N8496, N8497, N8500, N8501, N8502, N8503, N8504, N8505, N8506, N8507,
         N8508, N8509, N8510, N8511, N8512, N8513, N8514, N8515, N8516, N8517,
         N8518, N8519, N8522, N8525, N8528, N8531, N8534, N8537, N8538, N8539,
         N8540, N8541, N8545, N8546, N8547, N8548, N8551, N8552, N8553, N8554,
         N8555, N8558, N8561, N8564, N8565, N8566, N8569, N8572, N8575, N8578,
         N8579, N8580, N8583, N8586, N8589, N8592, N8595, N8598, N8601, N8604,
         N8607, N8608, N8609, N8610, N8615, N8616, N8617, N8618, N8619, N8624,
         N8625, N8626, N8627, N8632, N8633, N8634, N8637, N8638, N8639, N8644,
         N8645, N8646, N8647, N8648, N8653, N8654, N8655, N8660, N8663, N8666,
         N8669, N8672, N8675, N8678, N8681, N8684, N8687, N8690, N8693, N8696,
         N8699, N8702, N8705, N8708, N8711, N8714, N8717, N8718, N8721, N8724,
         N8727, N8730, N8733, N8734, N8735, N8738, N8741, N8744, N8747, N8750,
         N8753, N8754, N8755, N8756, N8757, N8760, N8763, N8766, N8769, N8772,
         N8775, N8778, N8781, N8784, N8787, N8790, N8793, N8796, N8799, N8802,
         N8805, N8808, N8811, N8814, N8815, N8816, N8817, N8818, N8840, N8857,
         N8861, N8862, N8863, N8864, N8865, N8866, N8871, N8874, N8878, N8879,
         N8880, N8881, N8882, N8883, N8884, N8885, N8886, N8887, N8888, N8898,
         N8902, N8920, N8924, N8927, N8931, N8943, N8950, N8956, N8959, N8960,
         N8963, N8966, N8991, N8992, N8995, N8996, N9001, N9005, N9024, N9025,
         N9029, N9035, N9053, N9054, N9064, N9065, N9066, N9067, N9068, N9071,
         N9072, N9073, N9074, N9077, N9079, N9082, N9083, N9086, N9087, N9088,
         N9089, N9092, N9093, N9094, N9095, N9098, N9099, N9103, N9107, N9111,
         N9117, N9127, N9146, N9149, N9159, N9160, N9161, N9165, N9169, N9173,
         N9179, N9180, N9181, N9182, N9183, N9193, N9203, N9206, N9220, N9223,
         N9234, N9235, N9236, N9237, N9238, N9242, N9243, N9244, N9245, N9246,
         N9247, N9248, N9249, N9250, N9251, N9252, N9256, N9257, N9258, N9259,
         N9260, N9261, N9262, N9265, N9268, N9271, N9272, N9273, N9274, N9275,
         N9276, N9280, N9285, N9286, N9287, N9288, N9290, N9292, N9294, N9296,
         N9297, N9298, N9299, N9300, N9301, N9307, N9314, N9315, N9318, N9319,
         N9320, N9321, N9322, N9323, N9324, N9326, N9332, N9339, N9344, N9352,
         N9354, N9356, N9358, N9359, N9360, N9361, N9362, N9363, N9364, N9365,
         N9366, N9367, N9368, N9369, N9370, N9371, N9372, N9375, N9381, N9382,
         N9383, N9384, N9385, N9392, N9393, N9394, N9395, N9396, N9397, N9398,
         N9399, N9400, N9401, N9402, N9407, N9408, N9412, N9413, N9414, N9415,
         N9416, N9417, N9418, N9419, N9420, N9421, N9422, N9423, N9426, N9429,
         N9432, N9435, N9442, N9445, N9454, N9455, N9456, N9459, N9460, N9461,
         N9462, N9465, N9466, N9467, N9468, N9473, N9476, N9477, N9478, N9485,
         N9488, N9493, N9494, N9495, N9498, N9499, N9500, N9505, N9506, N9507,
         N9508, N9509, N9514, N9515, N9516, N9517, N9520, N9526, N9531, N9539,
         N9540, N9541, N9543, N9551, N9555, N9556, N9557, N9560, N9561, N9562,
         N9563, N9564, N9565, N9566, N9567, N9568, N9569, N9570, N9571, N9575,
         N9579, N9581, N9582, N9585, N9591, N9592, N9593, N9594, N9595, N9596,
         N9597, N9598, N9599, N9600, N9601, N9602, N9603, N9604, N9605, N9608,
         N9611, N9612, N9613, N9614, N9615, N9616, N9617, N9618, N9621, N9622,
         N9623, N9624, N9626, N9629, N9632, N9635, N9642, N9645, N9646, N9649,
         N9650, N9653, N9656, N9659, N9660, N9661, N9662, N9663, N9666, N9667,
         N9670, N9671, N9674, N9675, N9678, N9679, N9682, N9685, N9690, N9691,
         N9692, N9695, N9698, N9702, N9707, N9710, N9711, N9714, N9715, N9716,
         N9717, N9720, N9721, N9722, N9723, N9726, N9727, N9732, N9733, N9734,
         N9735, N9736, N9737, N9738, N9739, N9740, N9741, N9742, N9754, N9758,
         N9762, N9763, N9764, N9765, N9766, N9767, N9768, N9769, N9773, N9774,
         N9775, N9779, N9784, N9785, N9786, N9790, N9791, N9795, N9796, N9797,
         N9798, N9799, N9800, N9801, N9802, N9803, N9805, N9806, N9809, N9813,
         N9814, N9815, N9816, N9817, N9820, N9825, N9826, N9827, N9828, N9829,
         N9830, N9835, N9836, N9837, N9838, N9846, N9847, N9862, N9863, N9866,
         N9873, N9876, N9890, N9891, N9892, N9893, N9894, N9895, N9896, N9897,
         N9898, N9899, N9900, N9901, N9902, N9903, N9904, N9905, N9906, N9907,
         N9908, N9909, N9910, N9911, N9917, N9923, N9924, N9925, N9932, N9935,
         N9938, N9939, N9945, N9946, N9947, N9948, N9949, N9953, N9954, N9955,
         N9956, N9957, N9958, N9959, N9960, N9961, N9964, N9967, N9968, N9969,
         N9970, N9971, N9972, N9973, N9974, N9975, N9976, N9977, N9978, N9979,
         N9982, N9983, N9986, N9989, N9992, N9995, N9996, N9997, N9998, N9999,
         N10002, N10003, N10006, N10007, N10010, N10013, N10014, N10015,
         N10016, N10017, N10018, N10019, N10020, N10021, N10022, N10023,
         N10024, N10026, N10028, N10032, N10033, N10034, N10035, N10036,
         N10037, N10038, N10039, N10040, N10041, N10042, N10043, N10050,
         N10053, N10054, N10055, N10056, N10057, N10058, N10059, N10060,
         N10061, N10062, N10067, N10070, N10073, N10076, N10077, N10082,
         N10083, N10084, N10085, N10086, N10093, N10094, N10105, N10106,
         N10107, N10108, N10113, N10114, N10115, N10116, N10119, N10124,
         N10130, N10131, N10132, N10133, N10134, N10135, N10136, N10137,
         N10138, N10139, N10140, N10141, N10148, N10155, N10156, N10157,
         N10158, N10159, N10160, N10161, N10162, N10163, N10164, N10165,
         N10170, N10173, N10176, N10177, N10178, N10179, N10180, N10183,
         N10186, N10189, N10192, N10195, N10196, N10197, N10200, N10203,
         N10204, N10205, N10206, N10212, N10213, N10230, N10231, N10232,
         N10233, N10234, N10237, N10238, N10239, N10240, N10241, N10242,
         N10247, N10248, N10259, N10264, N10265, N10266, N10267, N10268,
         N10269, N10270, N10271, N10272, N10273, N10278, N10279, N10280,
         N10281, N10282, N10283, N10287, N10288, N10289, N10290, N10291,
         N10292, N10293, N10294, N10295, N10296, N10299, N10300, N10301,
         N10306, N10307, N10308, N10311, N10314, N10315, N10316, N10317,
         N10318, N10321, N10324, N10325, N10326, N10327, N10328, N10329,
         N10330, N10331, N10332, N10333, N10334, N10337, N10338, N10339,
         N10340, N10341, N10344, N10354, N10357, N10360, N10367, N10375,
         N10381, N10388, N10391, N10399, N10402, N10406, N10409, N10412,
         N10415, N10419, N10422, N10425, N10428, N10431, N10432, N10437,
         N10438, N10439, N10440, N10441, N10444, N10445, N10450, N10451,
         N10455, N10456, N10465, N10466, N10479, N10497, N10509, N10512,
         N10515, N10516, N10517, N10518, N10519, N10522, N10525, N10528,
         N10531, N10534, N10535, N10536, N10539, N10542, N10543, N10544,
         N10545, N10546, N10547, N10548, N10549, N10550, N10551, N10552,
         N10553, N10554, N10555, N10556, N10557, N10558, N10559, N10560,
         N10561, N10562, N10563, N10564, N10565, N10566, N10567, N10568,
         N10569, N10570, N10571, N10572, N10573, N10577, N10581, N10582,
         N10583, N10587, N10588, N10589, N10594, N10595, N10596, N10597,
         N10598, N10602, N10609, N10610, N10621, N10626, N10627, N10629,
         N10631, N10637, N10638, N10639, N10640, N10642, N10643, N10644,
         N10645, N10647, N10648, N10649, N10652, N10659, N10662, N10665,
         N10668, N10671, N10672, N10673, N10674, N10675, N10678, N10681,
         N10682, N10683, N10684, N10685, N10686, N10687, N10688, N10689,
         N10690, N10691, N10694, N10695, N10696, N10697, N10698, N10701,
         N10705, N10707, N10708, N10709, N10710, N10719, N10720, N10730,
         N10731, N10737, N10738, N10739, N10746, N10747, N10748, N10749,
         N10750, N10753, N10754, N10764, N10765, N10766, N10767, N10768,
         N10769, N10770, N10771, N10772, N10773, N10774, N10775, N10776,
         N10778, N10781, N10784, N10789, N10792, N10796, N10797, N10798,
         N10799, N10800, N10803, N10806, N10809, N10812, N10815, N10816,
         N10817, N10820, N10823, N10824, N10825, N10826, N10832, N10833,
         N10834, N10835, N10836, N10845, N10846, N10857, N10862, N10863,
         N10864, N10865, N10866, N10867, N10872, N10873, N10874, N10875,
         N10876, N10879, N10882, N10883, N10884, N10885, N10886, N10887,
         N10888, N10889, N10890, N10891, N10892, N10895, N10896, N10897,
         N10898, N10899, N10902, N10909, N10910, N10915, N10916, N10917,
         N10918, N10919, N10922, N10923, N10928, N10931, N10934, N10935,
         N10936, N10937, N10938, N10941, N10944, N10947, N10950, N10953,
         N10954, N10955, N10958, N10961, N10962, N10963, N10964, N10969,
         N10970, N10981, N10986, N10987, N10988, N10989, N10990, N10991,
         N10992, N10995, N10998, N10999, N11000, N11001, N11002, N11003,
         N11004, N11005, N11006, N11007, N11008, N11011, N11012, N11013,
         N11014, N11015, N11018, N11023, N11024, N11027, N11028, N11029,
         N11030, N11031, N11034, N11035, N11040, N11041, N11042, N11043,
         N11044, N11047, N11050, N11053, N11056, N11059, N11062, N11065,
         N11066, N11067, N11070, N11073, N11074, N11075, N11076, N11077,
         N11078, N11095, N11098, N11099, N11100, N11103, N11106, N11107,
         N11108, N11109, N11110, N11111, N11112, N11113, N11114, N11115,
         N11116, N11117, N11118, N11119, N11120, N11121, N11122, N11123,
         N11124, N11127, N11130, N11137, N11138, N11139, N11140, N11141,
         N11142, N11143, N11144, N11145, N11152, N11153, N11154, N11155,
         N11156, N11159, N11162, N11165, N11168, N11171, N11174, N11177,
         N11180, N11183, N11184, N11185, N11186, N11187, N11188, N11205,
         N11210, N11211, N11212, N11213, N11214, N11215, N11216, N11217,
         N11218, N11219, N11220, N11222, N11223, N11224, N11225, N11226,
         N11227, N11228, N11229, N11231, N11232, N11233, N11236, N11239,
         N11242, N11243, N11244, N11245, N11246, N11250, N11252, N11257,
         N11260, N11261, N11262, N11263, N11264, N11265, N11267, N11268,
         N11269, N11270, N11272, N11277, N11278, N11279, N11280, N11282,
         N11283, N11284, N11285, N11286, N11288, N11289, N11290, N11291,
         N11292, N11293, N11294, N11295, N11296, N11297, N11298, N11299,
         N11302, N11307, N11308, N11309, N11312, N11313, N11314, N11315,
         N11316, N11317, N11320, N11321, N11323, N11327, N11328, N11329,
         N11331, N11335, N11336, N11337, N11338, N11339, N11341, N494_1,
         N494_2, N528_1, N528_2, N575_1, N575_2, N578_1, N578_2, N4303_1,
         N6762_1, N6762_2, N6762_3, N6767_1, N6768_1, N6768_2, N6769_1,
         N6769_2, N6769_3, N6771_1, N6772_1, N6772_2, N6773_1, N6773_2,
         N6775_1, N6776_1, N6776_2, N6778_1, N6779_1, N6781_1, N6784_1,
         N6784_2, N6784_3, N6788_1, N6789_1, N6789_2, N6790_1, N6790_2,
         N6790_3, N6792_1, N6793_1, N6793_2, N6795_1, N6833_1, N6833_2,
         N6837_1, N6838_1, N6838_2, N6840_1, N6841_1, N6843_1, N6845_1,
         N6845_2, N6845_3, N6849_1, N6850_1, N6850_2, N6851_1, N6851_2,
         N6851_3, N6853_1, N6854_1, N6854_2, N6855_1, N6855_2, N6857_1,
         N6858_1, N6858_2, N6860_1, N6861_1, N6863_1, N6867_1, N6867_2,
         N6871_1, N6872_1, N6872_2, N6874_1, N6875_1, N6877_1, N6881_1,
         N6881_2, N6881_3, N6885_1, N6886_1, N6886_2, N6887_1, N6887_2,
         N6887_3, N6889_1, N6890_1, N6890_2, N6892_1, N7057_1, N7057_2,
         N7061_1, N7062_1, N7062_2, N7063_1, N7063_2, N7063_3, N7065_1,
         N7066_1, N7066_2, N7067_1, N7067_2, N7067_3, N7100_1, N7100_2,
         N7100_3, N7104_1, N7105_1, N7105_2, N7106_1, N7106_2, N7106_3,
         N7609_1, N7609_2, N7609_3, N7620_1, N7620_2, N7620_3, N7649_1,
         N7649_2, N7655_1, N7655_2, N7655_3, N7668_1, N7668_2, N7671_1,
         N7671_2, N7671_3, N7825_1, N7825_2, N7826_1, N7826_2, N7826_3,
         N7852_1, N7852_2, N7852_3, N8114_1, N8114_2, N8117_1, N8117_2,
         N8117_3, N8134_1, N8134_2, N8146_1, N8146_2, N8166_1, N8166_2,
         N8169_1, N8169_2, N8169_3, N8186_1, N8186_2, N8196_1, N8196_2,
         N8204_1, N8280_1, N8281_1, N8282_1, N8283_1, N8284_1, N8285_1,
         N8333_1, N8333_2, N8338_1, N8339_1, N8339_2, N8341_1, N8342_1,
         N8344_1, N8349_1, N8350_1, N8350_2, N8351_1, N8351_2, N8351_3,
         N8353_1, N8354_1, N8354_2, N8356_1, N8365_1, N8365_2, N8370_1,
         N8371_1, N8371_2, N8373_1, N8374_1, N8376_1, N8379_1, N8380_1,
         N8380_2, N8381_1, N8381_2, N8381_3, N8383_1, N8384_1, N8384_2,
         N8386_1, N8387_1, N8387_2, N8389_1, N8391_1, N8405_1, N8405_2,
         N8410_1, N8411_1, N8411_2, N8412_1, N8412_2, N8412_3, N8416_1,
         N8417_1, N8417_2, N8418_1, N8418_2, N8418_3, N8430_1, N8430_2,
         N8434_1, N8435_1, N8435_2, N8437_1, N8438_1, N8440_1, N8444_1,
         N8444_2, N8444_3, N8448_1, N8449_1, N8449_2, N8450_1, N8450_2,
         N8450_3, N8452_1, N8453_1, N8453_2, N8455_1, N8483_1, N8484_1,
         N8485_1, N8485_2, N8489_1, N8490_1, N8490_2, N8492_1, N8493_1,
         N8495_1, N8497_1, N8497_2, N8497_3, N8501_1, N8502_1, N8502_2,
         N8503_1, N8503_2, N8503_3, N8505_1, N8506_1, N8506_2, N8507_1,
         N8507_2, N8509_1, N8510_1, N8510_2, N8512_1, N8513_1, N8515_1,
         N8539_1, N8540_1, N8541_1, N8541_2, N8546_1, N8547_1, N8547_2,
         N8548_1, N8548_2, N8548_3, N8552_1, N8553_1, N8553_2, N8554_1,
         N8554_2, N8554_3, N8578_1, N8579_1, N8861_1, N8862_1, N8863_1,
         N8864_1, N8865_1, N8866_1, N8898_1, N8898_2, N8902_1, N8902_2,
         N8902_3, N8920_1, N8920_2, N8927_1, N8927_2, N8927_3, N8950_1,
         N8950_2, N8956_1, N8956_2, N8956_3, N8963_1, N8963_2, N8966_1,
         N8966_2, N8966_3, N8991_1, N8992_1, N8995_1, N8995_2, N9001_1,
         N9001_2, N9001_3, N9024_1, N9025_1, N9029_1, N9029_2, N9035_1,
         N9035_2, N9035_3, N9053_1, N9054_1, N9099_1, N9099_2, N9107_1,
         N9117_1, N9117_2, N9149_1, N9149_2, N9161_1, N9161_2, N9169_1,
         N9183_1, N9183_2, N9203_1, N9203_2, N9206_1, N9206_2, N9206_3,
         N9223_1, N9223_2, N9280_1, N9280_2, N9280_3, N9285_1, N9285_2,
         N9285_3, N9286_1, N9286_2, N9287_1, N9307_1, N9307_2, N9307_3,
         N9314_1, N9314_2, N9315_1, N9369_1, N9370_1, N9371_1, N9372_1,
         N9396_1, N9397_1, N9398_1, N9399_1, N9419_1, N9420_1, N9421_1,
         N9422_1, N9602_1, N9603_1, N9604_1, N9605_1, N9612_1, N9613_1,
         N9614_1, N9615_1, N9621_1, N9622_1, N9623_1, N9624_1, N9626_1,
         N9626_2, N9626_3, N9629_1, N9629_2, N9632_1, N9679_1, N9679_2,
         N9685_1, N9685_2, N9685_3, N9734_1, N9734_2, N9734_3, N9735_1,
         N9735_2, N9735_3, N9790_1, N9790_2, N10013_1, N10014_1, N10014_2,
         N10015_1, N10015_2, N10015_3, N10016_1, N10017_1, N10017_2, N10018_1,
         N10019_1, N10019_2, N10020_1, N10021_1, N10021_2, N10022_1, N10022_2,
         N10022_3, N10040_1, N10041_1, N10041_2, N10043_1, N10056_1, N10058_1,
         N10059_1, N10059_2, N10061_1, N10101_1, N10101_2, N10101_3, N10102_1,
         N10102_2, N10102_3, N10103_1, N10103_2, N10103_3, N10104_1, N10104_2,
         N10104_3, N10116_1, N10116_2, N10119_1, N10140_1, N10140_2, N10141_1,
         N10141_2, N10148_1, N10278_1, N10278_2, N10278_3, N10279_1, N10279_2,
         N10280_1, N10287_1, N10287_2, N10287_3, N10288_1, N10288_2, N10289_1,
         N10388_1, N10388_2, N10399_1, N10399_2, N10402_1, N10402_2, N10406_1,
         N10406_2, N10406_3, N10409_1, N10409_2, N10412_1, N10419_1, N10419_2,
         N10419_3, N10422_1, N10422_2, N10425_1, N10577_1, N10581_1, N10582_1,
         N10594_1, N10594_2, N10594_3, N10595_1, N10595_2, N10596_1, N10647_1,
         N10648_1, N10649_1, N10659_1, N10659_2, N10659_3, N10662_1, N10662_2,
         N10665_1, N10739_1, N10739_2, N11152_1, N11153_1, N11154_1, N11155_1,
         N11205_1, N11205_2, N11222_1, N11223_1, N11224_1, N11225_1, N11226_1,
         N11227_1, N11228_1, N11229_1, N11252_1, N11252_2, N11257_1, N11257_2;

  BUFX2 gate1 ( .A(N1), .Y(N387) );
  BUFX2 gate2 ( .A(N1), .Y(N388) );
  INVX1 gate3 ( .A(N57), .Y(N467) );
  AND2X1 gate4 ( .A(N134), .B(N133), .Y(N469) );
  BUFX2 gate5 ( .A(N248), .Y(N478) );
  BUFX2 gate6 ( .A(N254), .Y(N482) );
  BUFX2 gate7 ( .A(N257), .Y(N484) );
  BUFX2 gate8 ( .A(N260), .Y(N486) );
  BUFX2 gate9 ( .A(N263), .Y(N489) );
  BUFX2 gate10 ( .A(N267), .Y(N492) );
  AND2X1 gate11_1 ( .A(N162), .B(N172), .Y(N494_1) );
  AND2X1 gate11_2 ( .A(N188), .B(N199), .Y(N494_2) );
  AND2X1 gate11 ( .A(N494_1), .B(N494_2), .Y(N494) );
  BUFX2 gate12 ( .A(N274), .Y(N501) );
  BUFX2 gate13 ( .A(N280), .Y(N505) );
  BUFX2 gate14 ( .A(N283), .Y(N507) );
  BUFX2 gate15 ( .A(N286), .Y(N509) );
  BUFX2 gate16 ( .A(N289), .Y(N511) );
  BUFX2 gate17 ( .A(N293), .Y(N513) );
  BUFX2 gate18 ( .A(N296), .Y(N515) );
  BUFX2 gate19 ( .A(N299), .Y(N517) );
  BUFX2 gate20 ( .A(N303), .Y(N519) );
  AND2X1 gate21_1 ( .A(N150), .B(N184), .Y(N528_1) );
  AND2X1 gate21_2 ( .A(N228), .B(N240), .Y(N528_2) );
  AND2X1 gate21 ( .A(N528_1), .B(N528_2), .Y(N528) );
  BUFX2 gate22 ( .A(N307), .Y(N535) );
  BUFX2 gate23 ( .A(N310), .Y(N537) );
  BUFX2 gate24 ( .A(N313), .Y(N539) );
  BUFX2 gate25 ( .A(N316), .Y(N541) );
  BUFX2 gate26 ( .A(N319), .Y(N543) );
  BUFX2 gate27 ( .A(N322), .Y(N545) );
  BUFX2 gate28 ( .A(N325), .Y(N547) );
  BUFX2 gate29 ( .A(N328), .Y(N549) );
  BUFX2 gate30 ( .A(N331), .Y(N551) );
  BUFX2 gate31 ( .A(N334), .Y(N553) );
  BUFX2 gate32 ( .A(N337), .Y(N556) );
  BUFX2 gate33 ( .A(N343), .Y(N559) );
  BUFX2 gate34 ( .A(N346), .Y(N561) );
  BUFX2 gate35 ( .A(N349), .Y(N563) );
  BUFX2 gate36 ( .A(N352), .Y(N565) );
  BUFX2 gate37 ( .A(N355), .Y(N567) );
  BUFX2 gate38 ( .A(N358), .Y(N569) );
  BUFX2 gate39 ( .A(N361), .Y(N571) );
  BUFX2 gate40 ( .A(N364), .Y(N573) );
  AND2X1 gate41_1 ( .A(N183), .B(N182), .Y(N575_1) );
  AND2X1 gate41_2 ( .A(N185), .B(N186), .Y(N575_2) );
  AND2X1 gate41 ( .A(N575_1), .B(N575_2), .Y(N575) );
  AND2X1 gate42_1 ( .A(N210), .B(N152), .Y(N578_1) );
  AND2X1 gate42_2 ( .A(N218), .B(N230), .Y(N578_2) );
  AND2X1 gate42 ( .A(N578_1), .B(N578_2), .Y(N578) );
  INVX1 gate43 ( .A(N15), .Y(N582) );
  INVX1 gate44 ( .A(N5), .Y(N585) );
  BUFX2 gate45 ( .A(N1), .Y(N590) );
  INVX1 gate46 ( .A(N5), .Y(N593) );
  INVX1 gate47 ( .A(N5), .Y(N596) );
  INVX1 gate48 ( .A(N289), .Y(N599) );
  INVX1 gate49 ( .A(N299), .Y(N604) );
  INVX1 gate50 ( .A(N303), .Y(N609) );
  BUFX2 gate51 ( .A(N38), .Y(N614) );
  BUFX2 gate52 ( .A(N15), .Y(N625) );
  NAND2X1 gate53 ( .A(N12), .B(N9), .Y(N628) );
  NAND2X1 gate54 ( .A(N12), .B(N9), .Y(N632) );
  BUFX2 gate55 ( .A(N38), .Y(N636) );
  INVX1 gate56 ( .A(N245), .Y(N641) );
  INVX1 gate57 ( .A(N248), .Y(N642) );
  BUFX2 gate58 ( .A(N251), .Y(N643) );
  INVX1 gate59 ( .A(N251), .Y(N644) );
  INVX1 gate60 ( .A(N254), .Y(N651) );
  BUFX2 gate61 ( .A(N106), .Y(N657) );
  INVX1 gate62 ( .A(N257), .Y(N660) );
  INVX1 gate63 ( .A(N260), .Y(N666) );
  INVX1 gate64 ( .A(N263), .Y(N672) );
  INVX1 gate65 ( .A(N267), .Y(N673) );
  INVX1 gate66 ( .A(N106), .Y(N674) );
  BUFX2 gate67 ( .A(N18), .Y(N676) );
  BUFX2 gate68 ( .A(N18), .Y(N682) );
  AND2X1 gate69 ( .A(N382), .B(N263), .Y(N688) );
  BUFX2 gate70 ( .A(N18), .Y(N689) );
  INVX1 gate71 ( .A(N18), .Y(N695) );
  NAND2X1 gate72 ( .A(N382), .B(N267), .Y(N700) );
  INVX1 gate73 ( .A(N271), .Y(N705) );
  INVX1 gate74 ( .A(N274), .Y(N706) );
  BUFX2 gate75 ( .A(N277), .Y(N707) );
  INVX1 gate76 ( .A(N277), .Y(N708) );
  INVX1 gate77 ( .A(N280), .Y(N715) );
  INVX1 gate78 ( .A(N283), .Y(N721) );
  INVX1 gate79 ( .A(N286), .Y(N727) );
  INVX1 gate80 ( .A(N289), .Y(N733) );
  INVX1 gate81 ( .A(N293), .Y(N734) );
  INVX1 gate82 ( .A(N296), .Y(N742) );
  INVX1 gate83 ( .A(N299), .Y(N748) );
  INVX1 gate84 ( .A(N303), .Y(N749) );
  BUFX2 gate85 ( .A(N367), .Y(N750) );
  INVX1 gate86 ( .A(N307), .Y(N758) );
  INVX1 gate87 ( .A(N310), .Y(N759) );
  INVX1 gate88 ( .A(N313), .Y(N762) );
  INVX1 gate89 ( .A(N316), .Y(N768) );
  INVX1 gate90 ( .A(N319), .Y(N774) );
  INVX1 gate91 ( .A(N322), .Y(N780) );
  INVX1 gate92 ( .A(N325), .Y(N786) );
  INVX1 gate93 ( .A(N328), .Y(N794) );
  INVX1 gate94 ( .A(N331), .Y(N800) );
  INVX1 gate95 ( .A(N334), .Y(N806) );
  INVX1 gate96 ( .A(N337), .Y(N812) );
  BUFX2 gate97 ( .A(N340), .Y(N813) );
  INVX1 gate98 ( .A(N340), .Y(N814) );
  INVX1 gate99 ( .A(N343), .Y(N821) );
  INVX1 gate100 ( .A(N346), .Y(N827) );
  INVX1 gate101 ( .A(N349), .Y(N833) );
  INVX1 gate102 ( .A(N352), .Y(N839) );
  INVX1 gate103 ( .A(N355), .Y(N845) );
  INVX1 gate104 ( .A(N358), .Y(N853) );
  INVX1 gate105 ( .A(N361), .Y(N859) );
  INVX1 gate106 ( .A(N364), .Y(N865) );
  BUFX2 gate107 ( .A(N367), .Y(N871) );
  NAND2X1 gate108 ( .A(N467), .B(N585), .Y(N881) );
  INVX1 gate109 ( .A(N528), .Y(N882) );
  INVX1 gate110 ( .A(N578), .Y(N883) );
  INVX1 gate111 ( .A(N575), .Y(N884) );
  INVX1 gate112 ( .A(N494), .Y(N885) );
  AND2X1 gate113 ( .A(N528), .B(N578), .Y(N886) );
  AND2X1 gate114 ( .A(N575), .B(N494), .Y(N887) );
  BUFX2 gate115 ( .A(N590), .Y(N889) );
  BUFX2 gate116 ( .A(N657), .Y(N945) );
  INVX1 gate117 ( .A(N688), .Y(N957) );
  AND2X1 gate118 ( .A(N382), .B(N641), .Y(N1028) );
  NAND2X1 gate119 ( .A(N382), .B(N705), .Y(N1029) );
  AND2X1 gate120 ( .A(N469), .B(N596), .Y(N1109) );
  NAND2X1 gate121 ( .A(N242), .B(N593), .Y(N1110) );
  INVX1 gate122 ( .A(N625), .Y(N1111) );
  NAND2X1 gate123 ( .A(N242), .B(N593), .Y(N1112) );
  NAND2X1 gate124 ( .A(N469), .B(N596), .Y(N1113) );
  INVX1 gate125 ( .A(N625), .Y(N1114) );
  INVX1 gate126 ( .A(N871), .Y(N1115) );
  BUFX2 gate127 ( .A(N590), .Y(N1116) );
  BUFX2 gate128 ( .A(N628), .Y(N1119) );
  BUFX2 gate129 ( .A(N682), .Y(N1125) );
  BUFX2 gate130 ( .A(N628), .Y(N1132) );
  BUFX2 gate131 ( .A(N682), .Y(N1136) );
  BUFX2 gate132 ( .A(N628), .Y(N1141) );
  BUFX2 gate133 ( .A(N682), .Y(N1147) );
  BUFX2 gate134 ( .A(N632), .Y(N1154) );
  BUFX2 gate135 ( .A(N676), .Y(N1160) );
  AND2X1 gate136 ( .A(N700), .B(N614), .Y(N1167) );
  AND2X1 gate137 ( .A(N700), .B(N614), .Y(N1174) );
  BUFX2 gate138 ( .A(N682), .Y(N1175) );
  BUFX2 gate139 ( .A(N676), .Y(N1182) );
  INVX1 gate140 ( .A(N657), .Y(N1189) );
  INVX1 gate141 ( .A(N676), .Y(N1194) );
  INVX1 gate142 ( .A(N682), .Y(N1199) );
  INVX1 gate143 ( .A(N689), .Y(N1206) );
  BUFX2 gate144 ( .A(N695), .Y(N1211) );
  INVX1 gate145 ( .A(N750), .Y(N1218) );
  INVX1 gate146 ( .A(N1028), .Y(N1222) );
  BUFX2 gate147 ( .A(N632), .Y(N1227) );
  BUFX2 gate148 ( .A(N676), .Y(N1233) );
  BUFX2 gate149 ( .A(N632), .Y(N1240) );
  BUFX2 gate150 ( .A(N676), .Y(N1244) );
  BUFX2 gate151 ( .A(N689), .Y(N1249) );
  BUFX2 gate152 ( .A(N689), .Y(N1256) );
  BUFX2 gate153 ( .A(N695), .Y(N1263) );
  BUFX2 gate154 ( .A(N689), .Y(N1270) );
  BUFX2 gate155 ( .A(N689), .Y(N1277) );
  BUFX2 gate156 ( .A(N700), .Y(N1284) );
  BUFX2 gate157 ( .A(N614), .Y(N1287) );
  BUFX2 gate158 ( .A(N666), .Y(N1290) );
  BUFX2 gate159 ( .A(N660), .Y(N1293) );
  BUFX2 gate160 ( .A(N651), .Y(N1296) );
  BUFX2 gate161 ( .A(N614), .Y(N1299) );
  BUFX2 gate162 ( .A(N644), .Y(N1302) );
  BUFX2 gate163 ( .A(N700), .Y(N1305) );
  BUFX2 gate164 ( .A(N614), .Y(N1308) );
  BUFX2 gate165 ( .A(N614), .Y(N1311) );
  BUFX2 gate166 ( .A(N666), .Y(N1314) );
  BUFX2 gate167 ( .A(N660), .Y(N1317) );
  BUFX2 gate168 ( .A(N651), .Y(N1320) );
  BUFX2 gate169 ( .A(N644), .Y(N1323) );
  BUFX2 gate170 ( .A(N609), .Y(N1326) );
  BUFX2 gate171 ( .A(N604), .Y(N1329) );
  BUFX2 gate172 ( .A(N742), .Y(N1332) );
  BUFX2 gate173 ( .A(N599), .Y(N1335) );
  BUFX2 gate174 ( .A(N727), .Y(N1338) );
  BUFX2 gate175 ( .A(N721), .Y(N1341) );
  BUFX2 gate176 ( .A(N715), .Y(N1344) );
  BUFX2 gate177 ( .A(N734), .Y(N1347) );
  BUFX2 gate178 ( .A(N708), .Y(N1350) );
  BUFX2 gate179 ( .A(N609), .Y(N1353) );
  BUFX2 gate180 ( .A(N604), .Y(N1356) );
  BUFX2 gate181 ( .A(N742), .Y(N1359) );
  BUFX2 gate182 ( .A(N734), .Y(N1362) );
  BUFX2 gate183 ( .A(N599), .Y(N1365) );
  BUFX2 gate184 ( .A(N727), .Y(N1368) );
  BUFX2 gate185 ( .A(N721), .Y(N1371) );
  BUFX2 gate186 ( .A(N715), .Y(N1374) );
  BUFX2 gate187 ( .A(N708), .Y(N1377) );
  BUFX2 gate188 ( .A(N806), .Y(N1380) );
  BUFX2 gate189 ( .A(N800), .Y(N1383) );
  BUFX2 gate190 ( .A(N794), .Y(N1386) );
  BUFX2 gate191 ( .A(N786), .Y(N1389) );
  BUFX2 gate192 ( .A(N780), .Y(N1392) );
  BUFX2 gate193 ( .A(N774), .Y(N1395) );
  BUFX2 gate194 ( .A(N768), .Y(N1398) );
  BUFX2 gate195 ( .A(N762), .Y(N1401) );
  BUFX2 gate196 ( .A(N806), .Y(N1404) );
  BUFX2 gate197 ( .A(N800), .Y(N1407) );
  BUFX2 gate198 ( .A(N794), .Y(N1410) );
  BUFX2 gate199 ( .A(N780), .Y(N1413) );
  BUFX2 gate200 ( .A(N774), .Y(N1416) );
  BUFX2 gate201 ( .A(N768), .Y(N1419) );
  BUFX2 gate202 ( .A(N762), .Y(N1422) );
  BUFX2 gate203 ( .A(N786), .Y(N1425) );
  BUFX2 gate204 ( .A(N636), .Y(N1428) );
  BUFX2 gate205 ( .A(N636), .Y(N1431) );
  BUFX2 gate206 ( .A(N865), .Y(N1434) );
  BUFX2 gate207 ( .A(N859), .Y(N1437) );
  BUFX2 gate208 ( .A(N853), .Y(N1440) );
  BUFX2 gate209 ( .A(N845), .Y(N1443) );
  BUFX2 gate210 ( .A(N839), .Y(N1446) );
  BUFX2 gate211 ( .A(N833), .Y(N1449) );
  BUFX2 gate212 ( .A(N827), .Y(N1452) );
  BUFX2 gate213 ( .A(N821), .Y(N1455) );
  BUFX2 gate214 ( .A(N814), .Y(N1458) );
  BUFX2 gate215 ( .A(N865), .Y(N1461) );
  BUFX2 gate216 ( .A(N859), .Y(N1464) );
  BUFX2 gate217 ( .A(N853), .Y(N1467) );
  BUFX2 gate218 ( .A(N839), .Y(N1470) );
  BUFX2 gate219 ( .A(N833), .Y(N1473) );
  BUFX2 gate220 ( .A(N827), .Y(N1476) );
  BUFX2 gate221 ( .A(N821), .Y(N1479) );
  BUFX2 gate222 ( .A(N845), .Y(N1482) );
  BUFX2 gate223 ( .A(N814), .Y(N1485) );
  INVX1 gate224 ( .A(N1109), .Y(N1489) );
  BUFX2 gate225 ( .A(N1116), .Y(N1490) );
  AND2X1 gate226 ( .A(N957), .B(N614), .Y(N1537) );
  AND2X1 gate227 ( .A(N614), .B(N957), .Y(N1551) );
  AND2X1 gate228 ( .A(N1029), .B(N636), .Y(N1649) );
  BUFX2 gate229 ( .A(N957), .Y(N1703) );
  NOR2X1 gate230 ( .A(N957), .B(N614), .Y(N1708) );
  BUFX2 gate231 ( .A(N957), .Y(N1713) );
  NOR2X1 gate232 ( .A(N614), .B(N957), .Y(N1721) );
  BUFX2 gate233 ( .A(N1029), .Y(N1758) );
  AND2X1 gate234 ( .A(N163), .B(N1116), .Y(N1781) );
  AND2X1 gate235 ( .A(N170), .B(N1125), .Y(N1782) );
  INVX1 gate236 ( .A(N1125), .Y(N1783) );
  INVX1 gate237 ( .A(N1136), .Y(N1789) );
  AND2X1 gate238 ( .A(N169), .B(N1125), .Y(N1793) );
  AND2X1 gate239 ( .A(N168), .B(N1125), .Y(N1794) );
  AND2X1 gate240 ( .A(N167), .B(N1125), .Y(N1795) );
  AND2X1 gate241 ( .A(N166), .B(N1136), .Y(N1796) );
  AND2X1 gate242 ( .A(N165), .B(N1136), .Y(N1797) );
  AND2X1 gate243 ( .A(N164), .B(N1136), .Y(N1798) );
  INVX1 gate244 ( .A(N1147), .Y(N1799) );
  INVX1 gate245 ( .A(N1160), .Y(N1805) );
  AND2X1 gate246 ( .A(N177), .B(N1147), .Y(N1811) );
  AND2X1 gate247 ( .A(N176), .B(N1147), .Y(N1812) );
  AND2X1 gate248 ( .A(N175), .B(N1147), .Y(N1813) );
  AND2X1 gate249 ( .A(N174), .B(N1147), .Y(N1814) );
  AND2X1 gate250 ( .A(N173), .B(N1147), .Y(N1815) );
  AND2X1 gate251 ( .A(N157), .B(N1160), .Y(N1816) );
  AND2X1 gate252 ( .A(N156), .B(N1160), .Y(N1817) );
  AND2X1 gate253 ( .A(N155), .B(N1160), .Y(N1818) );
  AND2X1 gate254 ( .A(N154), .B(N1160), .Y(N1819) );
  AND2X1 gate255 ( .A(N153), .B(N1160), .Y(N1820) );
  INVX1 gate256 ( .A(N1284), .Y(N1821) );
  INVX1 gate257 ( .A(N1287), .Y(N1822) );
  INVX1 gate258 ( .A(N1290), .Y(N1828) );
  INVX1 gate259 ( .A(N1293), .Y(N1829) );
  INVX1 gate260 ( .A(N1296), .Y(N1830) );
  INVX1 gate261 ( .A(N1299), .Y(N1832) );
  INVX1 gate262 ( .A(N1302), .Y(N1833) );
  INVX1 gate263 ( .A(N1305), .Y(N1834) );
  INVX1 gate264 ( .A(N1308), .Y(N1835) );
  INVX1 gate265 ( .A(N1311), .Y(N1839) );
  INVX1 gate266 ( .A(N1314), .Y(N1840) );
  INVX1 gate267 ( .A(N1317), .Y(N1841) );
  INVX1 gate268 ( .A(N1320), .Y(N1842) );
  INVX1 gate269 ( .A(N1323), .Y(N1843) );
  INVX1 gate270 ( .A(N1175), .Y(N1845) );
  INVX1 gate271 ( .A(N1182), .Y(N1851) );
  AND2X1 gate272 ( .A(N181), .B(N1175), .Y(N1857) );
  AND2X1 gate273 ( .A(N171), .B(N1175), .Y(N1858) );
  AND2X1 gate274 ( .A(N180), .B(N1175), .Y(N1859) );
  AND2X1 gate275 ( .A(N179), .B(N1175), .Y(N1860) );
  AND2X1 gate276 ( .A(N178), .B(N1175), .Y(N1861) );
  AND2X1 gate277 ( .A(N161), .B(N1182), .Y(N1862) );
  AND2X1 gate278 ( .A(N151), .B(N1182), .Y(N1863) );
  AND2X1 gate279 ( .A(N160), .B(N1182), .Y(N1864) );
  AND2X1 gate280 ( .A(N159), .B(N1182), .Y(N1865) );
  AND2X1 gate281 ( .A(N158), .B(N1182), .Y(N1866) );
  INVX1 gate282 ( .A(N1326), .Y(N1867) );
  INVX1 gate283 ( .A(N1329), .Y(N1868) );
  INVX1 gate284 ( .A(N1332), .Y(N1869) );
  INVX1 gate285 ( .A(N1335), .Y(N1870) );
  INVX1 gate286 ( .A(N1338), .Y(N1871) );
  INVX1 gate287 ( .A(N1341), .Y(N1872) );
  INVX1 gate288 ( .A(N1344), .Y(N1873) );
  INVX1 gate289 ( .A(N1347), .Y(N1874) );
  INVX1 gate290 ( .A(N1350), .Y(N1875) );
  INVX1 gate291 ( .A(N1353), .Y(N1876) );
  INVX1 gate292 ( .A(N1356), .Y(N1877) );
  INVX1 gate293 ( .A(N1359), .Y(N1878) );
  INVX1 gate294 ( .A(N1362), .Y(N1879) );
  INVX1 gate295 ( .A(N1365), .Y(N1880) );
  INVX1 gate296 ( .A(N1368), .Y(N1881) );
  INVX1 gate297 ( .A(N1371), .Y(N1882) );
  INVX1 gate298 ( .A(N1374), .Y(N1883) );
  INVX1 gate299 ( .A(N1377), .Y(N1884) );
  BUFX2 gate300 ( .A(N1199), .Y(N1885) );
  BUFX2 gate301 ( .A(N1194), .Y(N1892) );
  BUFX2 gate302 ( .A(N1199), .Y(N1899) );
  BUFX2 gate303 ( .A(N1194), .Y(N1906) );
  INVX1 gate304 ( .A(N1211), .Y(N1913) );
  BUFX2 gate305 ( .A(N1194), .Y(N1919) );
  AND2X1 gate306 ( .A(N44), .B(N1211), .Y(N1926) );
  AND2X1 gate307 ( .A(N41), .B(N1211), .Y(N1927) );
  AND2X1 gate308 ( .A(N29), .B(N1211), .Y(N1928) );
  AND2X1 gate309 ( .A(N26), .B(N1211), .Y(N1929) );
  AND2X1 gate310 ( .A(N23), .B(N1211), .Y(N1930) );
  INVX1 gate311 ( .A(N1380), .Y(N1931) );
  INVX1 gate312 ( .A(N1383), .Y(N1932) );
  INVX1 gate313 ( .A(N1386), .Y(N1933) );
  INVX1 gate314 ( .A(N1389), .Y(N1934) );
  INVX1 gate315 ( .A(N1392), .Y(N1935) );
  INVX1 gate316 ( .A(N1395), .Y(N1936) );
  INVX1 gate317 ( .A(N1398), .Y(N1937) );
  INVX1 gate318 ( .A(N1401), .Y(N1938) );
  INVX1 gate319 ( .A(N1404), .Y(N1939) );
  INVX1 gate320 ( .A(N1407), .Y(N1940) );
  INVX1 gate321 ( .A(N1410), .Y(N1941) );
  INVX1 gate322 ( .A(N1413), .Y(N1942) );
  INVX1 gate323 ( .A(N1416), .Y(N1943) );
  INVX1 gate324 ( .A(N1419), .Y(N1944) );
  INVX1 gate325 ( .A(N1422), .Y(N1945) );
  INVX1 gate326 ( .A(N1425), .Y(N1946) );
  INVX1 gate327 ( .A(N1233), .Y(N1947) );
  INVX1 gate328 ( .A(N1244), .Y(N1953) );
  AND2X1 gate329 ( .A(N209), .B(N1233), .Y(N1957) );
  AND2X1 gate330 ( .A(N216), .B(N1233), .Y(N1958) );
  AND2X1 gate331 ( .A(N215), .B(N1233), .Y(N1959) );
  AND2X1 gate332 ( .A(N214), .B(N1233), .Y(N1960) );
  AND2X1 gate333 ( .A(N213), .B(N1244), .Y(N1961) );
  AND2X1 gate334 ( .A(N212), .B(N1244), .Y(N1962) );
  AND2X1 gate335 ( .A(N211), .B(N1244), .Y(N1963) );
  INVX1 gate336 ( .A(N1428), .Y(N1965) );
  AND2X1 gate337 ( .A(N1222), .B(N636), .Y(N1966) );
  INVX1 gate338 ( .A(N1431), .Y(N1967) );
  INVX1 gate339 ( .A(N1434), .Y(N1968) );
  INVX1 gate340 ( .A(N1437), .Y(N1969) );
  INVX1 gate341 ( .A(N1440), .Y(N1970) );
  INVX1 gate342 ( .A(N1443), .Y(N1971) );
  INVX1 gate343 ( .A(N1446), .Y(N1972) );
  INVX1 gate344 ( .A(N1449), .Y(N1973) );
  INVX1 gate345 ( .A(N1452), .Y(N1974) );
  INVX1 gate346 ( .A(N1455), .Y(N1975) );
  INVX1 gate347 ( .A(N1458), .Y(N1976) );
  INVX1 gate348 ( .A(N1249), .Y(N1977) );
  INVX1 gate349 ( .A(N1256), .Y(N1983) );
  AND2X1 gate350 ( .A(N642), .B(N1249), .Y(N1989) );
  AND2X1 gate351 ( .A(N644), .B(N1249), .Y(N1990) );
  AND2X1 gate352 ( .A(N651), .B(N1249), .Y(N1991) );
  AND2X1 gate353 ( .A(N674), .B(N1249), .Y(N1992) );
  AND2X1 gate354 ( .A(N660), .B(N1249), .Y(N1993) );
  AND2X1 gate355 ( .A(N666), .B(N1256), .Y(N1994) );
  AND2X1 gate356 ( .A(N672), .B(N1256), .Y(N1995) );
  AND2X1 gate357 ( .A(N673), .B(N1256), .Y(N1996) );
  INVX1 gate358 ( .A(N1263), .Y(N1997) );
  BUFX2 gate359 ( .A(N1194), .Y(N2003) );
  AND2X1 gate360 ( .A(N47), .B(N1263), .Y(N2010) );
  AND2X1 gate361 ( .A(N35), .B(N1263), .Y(N2011) );
  AND2X1 gate362 ( .A(N32), .B(N1263), .Y(N2012) );
  AND2X1 gate363 ( .A(N50), .B(N1263), .Y(N2013) );
  AND2X1 gate364 ( .A(N66), .B(N1263), .Y(N2014) );
  INVX1 gate365 ( .A(N1461), .Y(N2015) );
  INVX1 gate366 ( .A(N1464), .Y(N2016) );
  INVX1 gate367 ( .A(N1467), .Y(N2017) );
  INVX1 gate368 ( .A(N1470), .Y(N2018) );
  INVX1 gate369 ( .A(N1473), .Y(N2019) );
  INVX1 gate370 ( .A(N1476), .Y(N2020) );
  INVX1 gate371 ( .A(N1479), .Y(N2021) );
  INVX1 gate372 ( .A(N1482), .Y(N2022) );
  INVX1 gate373 ( .A(N1485), .Y(N2023) );
  BUFX2 gate374 ( .A(N1206), .Y(N2024) );
  BUFX2 gate375 ( .A(N1206), .Y(N2031) );
  BUFX2 gate376 ( .A(N1206), .Y(N2038) );
  BUFX2 gate377 ( .A(N1206), .Y(N2045) );
  INVX1 gate378 ( .A(N1270), .Y(N2052) );
  INVX1 gate379 ( .A(N1277), .Y(N2058) );
  AND2X1 gate380 ( .A(N706), .B(N1270), .Y(N2064) );
  AND2X1 gate381 ( .A(N708), .B(N1270), .Y(N2065) );
  AND2X1 gate382 ( .A(N715), .B(N1270), .Y(N2066) );
  AND2X1 gate383 ( .A(N721), .B(N1270), .Y(N2067) );
  AND2X1 gate384 ( .A(N727), .B(N1270), .Y(N2068) );
  AND2X1 gate385 ( .A(N733), .B(N1277), .Y(N2069) );
  AND2X1 gate386 ( .A(N734), .B(N1277), .Y(N2070) );
  AND2X1 gate387 ( .A(N742), .B(N1277), .Y(N2071) );
  AND2X1 gate388 ( .A(N748), .B(N1277), .Y(N2072) );
  AND2X1 gate389 ( .A(N749), .B(N1277), .Y(N2073) );
  BUFX2 gate390 ( .A(N1189), .Y(N2074) );
  BUFX2 gate391 ( .A(N1189), .Y(N2081) );
  BUFX2 gate392 ( .A(N1222), .Y(N2086) );
  NAND2X1 gate393 ( .A(N1287), .B(N1821), .Y(N2107) );
  NAND2X1 gate394 ( .A(N1284), .B(N1822), .Y(N2108) );
  INVX1 gate395 ( .A(N1703), .Y(N2110) );
  NAND2X1 gate396 ( .A(N1703), .B(N1832), .Y(N2111) );
  NAND2X1 gate397 ( .A(N1308), .B(N1834), .Y(N2112) );
  NAND2X1 gate398 ( .A(N1305), .B(N1835), .Y(N2113) );
  INVX1 gate399 ( .A(N1713), .Y(N2114) );
  NAND2X1 gate400 ( .A(N1713), .B(N1839), .Y(N2115) );
  INVX1 gate401 ( .A(N1721), .Y(N2117) );
  INVX1 gate402 ( .A(N1758), .Y(N2171) );
  NAND2X1 gate403 ( .A(N1758), .B(N1965), .Y(N2172) );
  INVX1 gate404 ( .A(N1708), .Y(N2230) );
  BUFX2 gate405 ( .A(N1537), .Y(N2231) );
  BUFX2 gate406 ( .A(N1551), .Y(N2235) );
  OR2X1 gate407 ( .A(N1783), .B(N1782), .Y(N2239) );
  OR2X1 gate408 ( .A(N1783), .B(N1125), .Y(N2240) );
  OR2X1 gate409 ( .A(N1783), .B(N1793), .Y(N2241) );
  OR2X1 gate410 ( .A(N1783), .B(N1794), .Y(N2242) );
  OR2X1 gate411 ( .A(N1783), .B(N1795), .Y(N2243) );
  OR2X1 gate412 ( .A(N1789), .B(N1796), .Y(N2244) );
  OR2X1 gate413 ( .A(N1789), .B(N1797), .Y(N2245) );
  OR2X1 gate414 ( .A(N1789), .B(N1798), .Y(N2246) );
  OR2X1 gate415 ( .A(N1799), .B(N1811), .Y(N2247) );
  OR2X1 gate416 ( .A(N1799), .B(N1812), .Y(N2248) );
  OR2X1 gate417 ( .A(N1799), .B(N1813), .Y(N2249) );
  OR2X1 gate418 ( .A(N1799), .B(N1814), .Y(N2250) );
  OR2X1 gate419 ( .A(N1799), .B(N1815), .Y(N2251) );
  OR2X1 gate420 ( .A(N1805), .B(N1816), .Y(N2252) );
  OR2X1 gate421 ( .A(N1805), .B(N1817), .Y(N2253) );
  OR2X1 gate422 ( .A(N1805), .B(N1818), .Y(N2254) );
  OR2X1 gate423 ( .A(N1805), .B(N1819), .Y(N2255) );
  OR2X1 gate424 ( .A(N1805), .B(N1820), .Y(N2256) );
  NAND2X1 gate425 ( .A(N2107), .B(N2108), .Y(N2257) );
  INVX1 gate426 ( .A(N2074), .Y(N2267) );
  NAND2X1 gate427 ( .A(N1299), .B(N2110), .Y(N2268) );
  NAND2X1 gate428 ( .A(N2112), .B(N2113), .Y(N2269) );
  NAND2X1 gate429 ( .A(N1311), .B(N2114), .Y(N2274) );
  INVX1 gate430 ( .A(N2081), .Y(N2275) );
  AND2X1 gate431 ( .A(N141), .B(N1845), .Y(N2277) );
  AND2X1 gate432 ( .A(N147), .B(N1845), .Y(N2278) );
  AND2X1 gate433 ( .A(N138), .B(N1845), .Y(N2279) );
  AND2X1 gate434 ( .A(N144), .B(N1845), .Y(N2280) );
  AND2X1 gate435 ( .A(N135), .B(N1845), .Y(N2281) );
  AND2X1 gate436 ( .A(N141), .B(N1851), .Y(N2282) );
  AND2X1 gate437 ( .A(N147), .B(N1851), .Y(N2283) );
  AND2X1 gate438 ( .A(N138), .B(N1851), .Y(N2284) );
  AND2X1 gate439 ( .A(N144), .B(N1851), .Y(N2285) );
  AND2X1 gate440 ( .A(N135), .B(N1851), .Y(N2286) );
  INVX1 gate441 ( .A(N1885), .Y(N2287) );
  INVX1 gate442 ( .A(N1892), .Y(N2293) );
  AND2X1 gate443 ( .A(N103), .B(N1885), .Y(N2299) );
  AND2X1 gate444 ( .A(N130), .B(N1885), .Y(N2300) );
  AND2X1 gate445 ( .A(N127), .B(N1885), .Y(N2301) );
  AND2X1 gate446 ( .A(N124), .B(N1885), .Y(N2302) );
  AND2X1 gate447 ( .A(N100), .B(N1885), .Y(N2303) );
  AND2X1 gate448 ( .A(N103), .B(N1892), .Y(N2304) );
  AND2X1 gate449 ( .A(N130), .B(N1892), .Y(N2305) );
  AND2X1 gate450 ( .A(N127), .B(N1892), .Y(N2306) );
  AND2X1 gate451 ( .A(N124), .B(N1892), .Y(N2307) );
  AND2X1 gate452 ( .A(N100), .B(N1892), .Y(N2308) );
  INVX1 gate453 ( .A(N1899), .Y(N2309) );
  INVX1 gate454 ( .A(N1906), .Y(N2315) );
  AND2X1 gate455 ( .A(N115), .B(N1899), .Y(N2321) );
  AND2X1 gate456 ( .A(N118), .B(N1899), .Y(N2322) );
  AND2X1 gate457 ( .A(N97), .B(N1899), .Y(N2323) );
  AND2X1 gate458 ( .A(N94), .B(N1899), .Y(N2324) );
  AND2X1 gate459 ( .A(N121), .B(N1899), .Y(N2325) );
  AND2X1 gate460 ( .A(N115), .B(N1906), .Y(N2326) );
  AND2X1 gate461 ( .A(N118), .B(N1906), .Y(N2327) );
  AND2X1 gate462 ( .A(N97), .B(N1906), .Y(N2328) );
  AND2X1 gate463 ( .A(N94), .B(N1906), .Y(N2329) );
  AND2X1 gate464 ( .A(N121), .B(N1906), .Y(N2330) );
  INVX1 gate465 ( .A(N1919), .Y(N2331) );
  AND2X1 gate466 ( .A(N208), .B(N1913), .Y(N2337) );
  AND2X1 gate467 ( .A(N198), .B(N1913), .Y(N2338) );
  AND2X1 gate468 ( .A(N207), .B(N1913), .Y(N2339) );
  AND2X1 gate469 ( .A(N206), .B(N1913), .Y(N2340) );
  AND2X1 gate470 ( .A(N205), .B(N1913), .Y(N2341) );
  AND2X1 gate471 ( .A(N44), .B(N1919), .Y(N2342) );
  AND2X1 gate472 ( .A(N41), .B(N1919), .Y(N2343) );
  AND2X1 gate473 ( .A(N29), .B(N1919), .Y(N2344) );
  AND2X1 gate474 ( .A(N26), .B(N1919), .Y(N2345) );
  AND2X1 gate475 ( .A(N23), .B(N1919), .Y(N2346) );
  OR2X1 gate476 ( .A(N1947), .B(N1233), .Y(N2347) );
  OR2X1 gate477 ( .A(N1947), .B(N1957), .Y(N2348) );
  OR2X1 gate478 ( .A(N1947), .B(N1958), .Y(N2349) );
  OR2X1 gate479 ( .A(N1947), .B(N1959), .Y(N2350) );
  OR2X1 gate480 ( .A(N1947), .B(N1960), .Y(N2351) );
  OR2X1 gate481 ( .A(N1953), .B(N1961), .Y(N2352) );
  OR2X1 gate482 ( .A(N1953), .B(N1962), .Y(N2353) );
  OR2X1 gate483 ( .A(N1953), .B(N1963), .Y(N2354) );
  NAND2X1 gate484 ( .A(N1428), .B(N2171), .Y(N2355) );
  INVX1 gate485 ( .A(N2086), .Y(N2356) );
  NAND2X1 gate486 ( .A(N2086), .B(N1967), .Y(N2357) );
  AND2X1 gate487 ( .A(N114), .B(N1977), .Y(N2358) );
  AND2X1 gate488 ( .A(N113), .B(N1977), .Y(N2359) );
  AND2X1 gate489 ( .A(N111), .B(N1977), .Y(N2360) );
  AND2X1 gate490 ( .A(N87), .B(N1977), .Y(N2361) );
  AND2X1 gate491 ( .A(N112), .B(N1977), .Y(N2362) );
  AND2X1 gate492 ( .A(N88), .B(N1983), .Y(N2363) );
  AND2X1 gate493 ( .A(N245), .B(N1983), .Y(N2364) );
  AND2X1 gate494 ( .A(N271), .B(N1983), .Y(N2365) );
  AND2X1 gate495 ( .A(N759), .B(N1983), .Y(N2366) );
  AND2X1 gate496 ( .A(N70), .B(N1983), .Y(N2367) );
  INVX1 gate497 ( .A(N2003), .Y(N2368) );
  AND2X1 gate498 ( .A(N193), .B(N1997), .Y(N2374) );
  AND2X1 gate499 ( .A(N192), .B(N1997), .Y(N2375) );
  AND2X1 gate500 ( .A(N191), .B(N1997), .Y(N2376) );
  AND2X1 gate501 ( .A(N190), .B(N1997), .Y(N2377) );
  AND2X1 gate502 ( .A(N189), .B(N1997), .Y(N2378) );
  AND2X1 gate503 ( .A(N47), .B(N2003), .Y(N2379) );
  AND2X1 gate504 ( .A(N35), .B(N2003), .Y(N2380) );
  AND2X1 gate505 ( .A(N32), .B(N2003), .Y(N2381) );
  AND2X1 gate506 ( .A(N50), .B(N2003), .Y(N2382) );
  AND2X1 gate507 ( .A(N66), .B(N2003), .Y(N2383) );
  INVX1 gate508 ( .A(N2024), .Y(N2384) );
  INVX1 gate509 ( .A(N2031), .Y(N2390) );
  AND2X1 gate510 ( .A(N58), .B(N2024), .Y(N2396) );
  AND2X1 gate511 ( .A(N77), .B(N2024), .Y(N2397) );
  AND2X1 gate512 ( .A(N78), .B(N2024), .Y(N2398) );
  AND2X1 gate513 ( .A(N59), .B(N2024), .Y(N2399) );
  AND2X1 gate514 ( .A(N81), .B(N2024), .Y(N2400) );
  AND2X1 gate515 ( .A(N80), .B(N2031), .Y(N2401) );
  AND2X1 gate516 ( .A(N79), .B(N2031), .Y(N2402) );
  AND2X1 gate517 ( .A(N60), .B(N2031), .Y(N2403) );
  AND2X1 gate518 ( .A(N61), .B(N2031), .Y(N2404) );
  AND2X1 gate519 ( .A(N62), .B(N2031), .Y(N2405) );
  INVX1 gate520 ( .A(N2038), .Y(N2406) );
  INVX1 gate521 ( .A(N2045), .Y(N2412) );
  AND2X1 gate522 ( .A(N69), .B(N2038), .Y(N2418) );
  AND2X1 gate523 ( .A(N70), .B(N2038), .Y(N2419) );
  AND2X1 gate524 ( .A(N74), .B(N2038), .Y(N2420) );
  AND2X1 gate525 ( .A(N76), .B(N2038), .Y(N2421) );
  AND2X1 gate526 ( .A(N75), .B(N2038), .Y(N2422) );
  AND2X1 gate527 ( .A(N73), .B(N2045), .Y(N2423) );
  AND2X1 gate528 ( .A(N53), .B(N2045), .Y(N2424) );
  AND2X1 gate529 ( .A(N54), .B(N2045), .Y(N2425) );
  AND2X1 gate530 ( .A(N55), .B(N2045), .Y(N2426) );
  AND2X1 gate531 ( .A(N56), .B(N2045), .Y(N2427) );
  AND2X1 gate532 ( .A(N82), .B(N2052), .Y(N2428) );
  AND2X1 gate533 ( .A(N65), .B(N2052), .Y(N2429) );
  AND2X1 gate534 ( .A(N83), .B(N2052), .Y(N2430) );
  AND2X1 gate535 ( .A(N84), .B(N2052), .Y(N2431) );
  AND2X1 gate536 ( .A(N85), .B(N2052), .Y(N2432) );
  AND2X1 gate537 ( .A(N64), .B(N2058), .Y(N2433) );
  AND2X1 gate538 ( .A(N63), .B(N2058), .Y(N2434) );
  AND2X1 gate539 ( .A(N86), .B(N2058), .Y(N2435) );
  AND2X1 gate540 ( .A(N109), .B(N2058), .Y(N2436) );
  AND2X1 gate541 ( .A(N110), .B(N2058), .Y(N2437) );
  AND2X1 gate542 ( .A(N2239), .B(N1119), .Y(N2441) );
  AND2X1 gate543 ( .A(N2240), .B(N1119), .Y(N2442) );
  AND2X1 gate544 ( .A(N2241), .B(N1119), .Y(N2446) );
  AND2X1 gate545 ( .A(N2242), .B(N1119), .Y(N2450) );
  AND2X1 gate546 ( .A(N2243), .B(N1119), .Y(N2454) );
  AND2X1 gate547 ( .A(N2244), .B(N1132), .Y(N2458) );
  AND2X1 gate548 ( .A(N2247), .B(N1141), .Y(N2462) );
  AND2X1 gate549 ( .A(N2248), .B(N1141), .Y(N2466) );
  AND2X1 gate550 ( .A(N2249), .B(N1141), .Y(N2470) );
  AND2X1 gate551 ( .A(N2250), .B(N1141), .Y(N2474) );
  AND2X1 gate552 ( .A(N2251), .B(N1141), .Y(N2478) );
  AND2X1 gate553 ( .A(N2252), .B(N1154), .Y(N2482) );
  AND2X1 gate554 ( .A(N2253), .B(N1154), .Y(N2488) );
  AND2X1 gate555 ( .A(N2254), .B(N1154), .Y(N2496) );
  AND2X1 gate556 ( .A(N2255), .B(N1154), .Y(N2502) );
  AND2X1 gate557 ( .A(N2256), .B(N1154), .Y(N2508) );
  NAND2X1 gate558 ( .A(N2268), .B(N2111), .Y(N2523) );
  NAND2X1 gate559 ( .A(N2274), .B(N2115), .Y(N2533) );
  INVX1 gate560 ( .A(N2235), .Y(N2537) );
  OR2X1 gate561 ( .A(N2278), .B(N1858), .Y(N2538) );
  OR2X1 gate562 ( .A(N2279), .B(N1859), .Y(N2542) );
  OR2X1 gate563 ( .A(N2280), .B(N1860), .Y(N2546) );
  OR2X1 gate564 ( .A(N2281), .B(N1861), .Y(N2550) );
  OR2X1 gate565 ( .A(N2283), .B(N1863), .Y(N2554) );
  OR2X1 gate566 ( .A(N2284), .B(N1864), .Y(N2561) );
  OR2X1 gate567 ( .A(N2285), .B(N1865), .Y(N2567) );
  OR2X1 gate568 ( .A(N2286), .B(N1866), .Y(N2573) );
  OR2X1 gate569 ( .A(N2338), .B(N1927), .Y(N2604) );
  OR2X1 gate570 ( .A(N2339), .B(N1928), .Y(N2607) );
  OR2X1 gate571 ( .A(N2340), .B(N1929), .Y(N2611) );
  OR2X1 gate572 ( .A(N2341), .B(N1930), .Y(N2615) );
  AND2X1 gate573 ( .A(N2348), .B(N1227), .Y(N2619) );
  AND2X1 gate574 ( .A(N2349), .B(N1227), .Y(N2626) );
  AND2X1 gate575 ( .A(N2350), .B(N1227), .Y(N2632) );
  AND2X1 gate576 ( .A(N2351), .B(N1227), .Y(N2638) );
  AND2X1 gate577 ( .A(N2352), .B(N1240), .Y(N2644) );
  NAND2X1 gate578 ( .A(N2355), .B(N2172), .Y(N2650) );
  NAND2X1 gate579 ( .A(N1431), .B(N2356), .Y(N2653) );
  OR2X1 gate580 ( .A(N2359), .B(N1990), .Y(N2654) );
  OR2X1 gate581 ( .A(N2360), .B(N1991), .Y(N2658) );
  OR2X1 gate582 ( .A(N2361), .B(N1992), .Y(N2662) );
  OR2X1 gate583 ( .A(N2362), .B(N1993), .Y(N2666) );
  OR2X1 gate584 ( .A(N2363), .B(N1994), .Y(N2670) );
  OR2X1 gate585 ( .A(N2366), .B(N1256), .Y(N2674) );
  OR2X1 gate586 ( .A(N2367), .B(N1256), .Y(N2680) );
  OR2X1 gate587 ( .A(N2374), .B(N2010), .Y(N2688) );
  OR2X1 gate588 ( .A(N2375), .B(N2011), .Y(N2692) );
  OR2X1 gate589 ( .A(N2376), .B(N2012), .Y(N2696) );
  OR2X1 gate590 ( .A(N2377), .B(N2013), .Y(N2700) );
  OR2X1 gate591 ( .A(N2378), .B(N2014), .Y(N2704) );
  AND2X1 gate592 ( .A(N2347), .B(N1227), .Y(N2728) );
  OR2X1 gate593 ( .A(N2429), .B(N2065), .Y(N2729) );
  OR2X1 gate594 ( .A(N2430), .B(N2066), .Y(N2733) );
  OR2X1 gate595 ( .A(N2431), .B(N2067), .Y(N2737) );
  OR2X1 gate596 ( .A(N2432), .B(N2068), .Y(N2741) );
  OR2X1 gate597 ( .A(N2433), .B(N2069), .Y(N2745) );
  OR2X1 gate598 ( .A(N2434), .B(N2070), .Y(N2749) );
  OR2X1 gate599 ( .A(N2435), .B(N2071), .Y(N2753) );
  OR2X1 gate600 ( .A(N2436), .B(N2072), .Y(N2757) );
  OR2X1 gate601 ( .A(N2437), .B(N2073), .Y(N2761) );
  INVX1 gate602 ( .A(N2231), .Y(N2765) );
  AND2X1 gate603 ( .A(N2354), .B(N1240), .Y(N2766) );
  AND2X1 gate604 ( .A(N2353), .B(N1240), .Y(N2769) );
  AND2X1 gate605 ( .A(N2246), .B(N1132), .Y(N2772) );
  AND2X1 gate606 ( .A(N2245), .B(N1132), .Y(N2775) );
  OR2X1 gate607 ( .A(N2282), .B(N1862), .Y(N2778) );
  OR2X1 gate608 ( .A(N2358), .B(N1989), .Y(N2781) );
  OR2X1 gate609 ( .A(N2365), .B(N1996), .Y(N2784) );
  OR2X1 gate610 ( .A(N2364), .B(N1995), .Y(N2787) );
  OR2X1 gate611 ( .A(N2337), .B(N1926), .Y(N2790) );
  OR2X1 gate612 ( .A(N2277), .B(N1857), .Y(N2793) );
  OR2X1 gate613 ( .A(N2428), .B(N2064), .Y(N2796) );
  AND2X1 gate614 ( .A(N2257), .B(N1537), .Y(N2866) );
  AND2X1 gate615 ( .A(N2257), .B(N1537), .Y(N2867) );
  AND2X1 gate616 ( .A(N2257), .B(N1537), .Y(N2868) );
  AND2X1 gate617 ( .A(N2257), .B(N1537), .Y(N2869) );
  AND2X1 gate618 ( .A(N2269), .B(N1551), .Y(N2878) );
  AND2X1 gate619 ( .A(N204), .B(N2287), .Y(N2913) );
  AND2X1 gate620 ( .A(N203), .B(N2287), .Y(N2914) );
  AND2X1 gate621 ( .A(N202), .B(N2287), .Y(N2915) );
  AND2X1 gate622 ( .A(N201), .B(N2287), .Y(N2916) );
  AND2X1 gate623 ( .A(N200), .B(N2287), .Y(N2917) );
  AND2X1 gate624 ( .A(N235), .B(N2293), .Y(N2918) );
  AND2X1 gate625 ( .A(N234), .B(N2293), .Y(N2919) );
  AND2X1 gate626 ( .A(N233), .B(N2293), .Y(N2920) );
  AND2X1 gate627 ( .A(N232), .B(N2293), .Y(N2921) );
  AND2X1 gate628 ( .A(N231), .B(N2293), .Y(N2922) );
  AND2X1 gate629 ( .A(N197), .B(N2309), .Y(N2923) );
  AND2X1 gate630 ( .A(N187), .B(N2309), .Y(N2924) );
  AND2X1 gate631 ( .A(N196), .B(N2309), .Y(N2925) );
  AND2X1 gate632 ( .A(N195), .B(N2309), .Y(N2926) );
  AND2X1 gate633 ( .A(N194), .B(N2309), .Y(N2927) );
  AND2X1 gate634 ( .A(N227), .B(N2315), .Y(N2928) );
  AND2X1 gate635 ( .A(N217), .B(N2315), .Y(N2929) );
  AND2X1 gate636 ( .A(N226), .B(N2315), .Y(N2930) );
  AND2X1 gate637 ( .A(N225), .B(N2315), .Y(N2931) );
  AND2X1 gate638 ( .A(N224), .B(N2315), .Y(N2932) );
  AND2X1 gate639 ( .A(N239), .B(N2331), .Y(N2933) );
  AND2X1 gate640 ( .A(N229), .B(N2331), .Y(N2934) );
  AND2X1 gate641 ( .A(N238), .B(N2331), .Y(N2935) );
  AND2X1 gate642 ( .A(N237), .B(N2331), .Y(N2936) );
  AND2X1 gate643 ( .A(N236), .B(N2331), .Y(N2937) );
  NAND2X1 gate644 ( .A(N2653), .B(N2357), .Y(N2988) );
  AND2X1 gate645 ( .A(N223), .B(N2368), .Y(N3005) );
  AND2X1 gate646 ( .A(N222), .B(N2368), .Y(N3006) );
  AND2X1 gate647 ( .A(N221), .B(N2368), .Y(N3007) );
  AND2X1 gate648 ( .A(N220), .B(N2368), .Y(N3008) );
  AND2X1 gate649 ( .A(N219), .B(N2368), .Y(N3009) );
  AND2X1 gate650 ( .A(N812), .B(N2384), .Y(N3020) );
  AND2X1 gate651 ( .A(N814), .B(N2384), .Y(N3021) );
  AND2X1 gate652 ( .A(N821), .B(N2384), .Y(N3022) );
  AND2X1 gate653 ( .A(N827), .B(N2384), .Y(N3023) );
  AND2X1 gate654 ( .A(N833), .B(N2384), .Y(N3024) );
  AND2X1 gate655 ( .A(N839), .B(N2390), .Y(N3025) );
  AND2X1 gate656 ( .A(N845), .B(N2390), .Y(N3026) );
  AND2X1 gate657 ( .A(N853), .B(N2390), .Y(N3027) );
  AND2X1 gate658 ( .A(N859), .B(N2390), .Y(N3028) );
  AND2X1 gate659 ( .A(N865), .B(N2390), .Y(N3029) );
  AND2X1 gate660 ( .A(N758), .B(N2406), .Y(N3032) );
  AND2X1 gate661 ( .A(N759), .B(N2406), .Y(N3033) );
  AND2X1 gate662 ( .A(N762), .B(N2406), .Y(N3034) );
  AND2X1 gate663 ( .A(N768), .B(N2406), .Y(N3035) );
  AND2X1 gate664 ( .A(N774), .B(N2406), .Y(N3036) );
  AND2X1 gate665 ( .A(N780), .B(N2412), .Y(N3037) );
  AND2X1 gate666 ( .A(N786), .B(N2412), .Y(N3038) );
  AND2X1 gate667 ( .A(N794), .B(N2412), .Y(N3039) );
  AND2X1 gate668 ( .A(N800), .B(N2412), .Y(N3040) );
  AND2X1 gate669 ( .A(N806), .B(N2412), .Y(N3041) );
  BUFX2 gate670 ( .A(N2257), .Y(N3061) );
  BUFX2 gate671 ( .A(N2257), .Y(N3064) );
  BUFX2 gate672 ( .A(N2269), .Y(N3067) );
  BUFX2 gate673 ( .A(N2269), .Y(N3070) );
  INVX1 gate674 ( .A(N2728), .Y(N3073) );
  INVX1 gate675 ( .A(N2441), .Y(N3080) );
  AND2X1 gate676 ( .A(N666), .B(N2644), .Y(N3096) );
  AND2X1 gate677 ( .A(N660), .B(N2638), .Y(N3097) );
  AND2X1 gate678 ( .A(N1189), .B(N2632), .Y(N3101) );
  AND2X1 gate679 ( .A(N651), .B(N2626), .Y(N3107) );
  AND2X1 gate680 ( .A(N644), .B(N2619), .Y(N3114) );
  AND2X1 gate681 ( .A(N2523), .B(N2257), .Y(N3122) );
  OR2X1 gate682 ( .A(N1167), .B(N2866), .Y(N3126) );
  AND2X1 gate683 ( .A(N2523), .B(N2257), .Y(N3130) );
  OR2X1 gate684 ( .A(N1167), .B(N2869), .Y(N3131) );
  AND2X1 gate685 ( .A(N2523), .B(N2257), .Y(N3134) );
  INVX1 gate686 ( .A(N2533), .Y(N3135) );
  AND2X1 gate687 ( .A(N666), .B(N2644), .Y(N3136) );
  AND2X1 gate688 ( .A(N660), .B(N2638), .Y(N3137) );
  AND2X1 gate689 ( .A(N1189), .B(N2632), .Y(N3140) );
  AND2X1 gate690 ( .A(N651), .B(N2626), .Y(N3144) );
  AND2X1 gate691 ( .A(N644), .B(N2619), .Y(N3149) );
  AND2X1 gate692 ( .A(N2533), .B(N2269), .Y(N3155) );
  OR2X1 gate693 ( .A(N1174), .B(N2878), .Y(N3159) );
  INVX1 gate694 ( .A(N2778), .Y(N3167) );
  AND2X1 gate695 ( .A(N609), .B(N2508), .Y(N3168) );
  AND2X1 gate696 ( .A(N604), .B(N2502), .Y(N3169) );
  AND2X1 gate697 ( .A(N742), .B(N2496), .Y(N3173) );
  AND2X1 gate698 ( .A(N734), .B(N2488), .Y(N3178) );
  AND2X1 gate699 ( .A(N599), .B(N2482), .Y(N3184) );
  AND2X1 gate700 ( .A(N727), .B(N2573), .Y(N3185) );
  AND2X1 gate701 ( .A(N721), .B(N2567), .Y(N3189) );
  AND2X1 gate702 ( .A(N715), .B(N2561), .Y(N3195) );
  AND2X1 gate703 ( .A(N708), .B(N2554), .Y(N3202) );
  AND2X1 gate704 ( .A(N609), .B(N2508), .Y(N3210) );
  AND2X1 gate705 ( .A(N604), .B(N2502), .Y(N3211) );
  AND2X1 gate706 ( .A(N742), .B(N2496), .Y(N3215) );
  AND2X1 gate707 ( .A(N2488), .B(N734), .Y(N3221) );
  AND2X1 gate708 ( .A(N599), .B(N2482), .Y(N3228) );
  AND2X1 gate709 ( .A(N727), .B(N2573), .Y(N3229) );
  AND2X1 gate710 ( .A(N721), .B(N2567), .Y(N3232) );
  AND2X1 gate711 ( .A(N715), .B(N2561), .Y(N3236) );
  AND2X1 gate712 ( .A(N708), .B(N2554), .Y(N3241) );
  OR2X1 gate713 ( .A(N2913), .B(N2299), .Y(N3247) );
  OR2X1 gate714 ( .A(N2914), .B(N2300), .Y(N3251) );
  OR2X1 gate715 ( .A(N2915), .B(N2301), .Y(N3255) );
  OR2X1 gate716 ( .A(N2916), .B(N2302), .Y(N3259) );
  OR2X1 gate717 ( .A(N2917), .B(N2303), .Y(N3263) );
  OR2X1 gate718 ( .A(N2918), .B(N2304), .Y(N3267) );
  OR2X1 gate719 ( .A(N2919), .B(N2305), .Y(N3273) );
  OR2X1 gate720 ( .A(N2920), .B(N2306), .Y(N3281) );
  OR2X1 gate721 ( .A(N2921), .B(N2307), .Y(N3287) );
  OR2X1 gate722 ( .A(N2922), .B(N2308), .Y(N3293) );
  OR2X1 gate723 ( .A(N2924), .B(N2322), .Y(N3299) );
  OR2X1 gate724 ( .A(N2925), .B(N2323), .Y(N3303) );
  OR2X1 gate725 ( .A(N2926), .B(N2324), .Y(N3307) );
  OR2X1 gate726 ( .A(N2927), .B(N2325), .Y(N3311) );
  OR2X1 gate727 ( .A(N2929), .B(N2327), .Y(N3315) );
  OR2X1 gate728 ( .A(N2930), .B(N2328), .Y(N3322) );
  OR2X1 gate729 ( .A(N2931), .B(N2329), .Y(N3328) );
  OR2X1 gate730 ( .A(N2932), .B(N2330), .Y(N3334) );
  OR2X1 gate731 ( .A(N2934), .B(N2343), .Y(N3340) );
  OR2X1 gate732 ( .A(N2935), .B(N2344), .Y(N3343) );
  OR2X1 gate733 ( .A(N2936), .B(N2345), .Y(N3349) );
  OR2X1 gate734 ( .A(N2937), .B(N2346), .Y(N3355) );
  AND2X1 gate735 ( .A(N2761), .B(N2478), .Y(N3361) );
  AND2X1 gate736 ( .A(N2757), .B(N2474), .Y(N3362) );
  AND2X1 gate737 ( .A(N2753), .B(N2470), .Y(N3363) );
  AND2X1 gate738 ( .A(N2749), .B(N2466), .Y(N3364) );
  AND2X1 gate739 ( .A(N2745), .B(N2462), .Y(N3365) );
  AND2X1 gate740 ( .A(N2741), .B(N2550), .Y(N3366) );
  AND2X1 gate741 ( .A(N2737), .B(N2546), .Y(N3367) );
  AND2X1 gate742 ( .A(N2733), .B(N2542), .Y(N3368) );
  AND2X1 gate743 ( .A(N2729), .B(N2538), .Y(N3369) );
  AND2X1 gate744 ( .A(N2670), .B(N2458), .Y(N3370) );
  AND2X1 gate745 ( .A(N2666), .B(N2454), .Y(N3371) );
  AND2X1 gate746 ( .A(N2662), .B(N2450), .Y(N3372) );
  AND2X1 gate747 ( .A(N2658), .B(N2446), .Y(N3373) );
  AND2X1 gate748 ( .A(N2654), .B(N2442), .Y(N3374) );
  AND2X1 gate749 ( .A(N2988), .B(N2650), .Y(N3375) );
  AND2X1 gate750 ( .A(N2650), .B(N1966), .Y(N3379) );
  INVX1 gate751 ( .A(N2781), .Y(N3380) );
  AND2X1 gate752 ( .A(N695), .B(N2604), .Y(N3381) );
  OR2X1 gate753 ( .A(N3005), .B(N2379), .Y(N3384) );
  OR2X1 gate754 ( .A(N3006), .B(N2380), .Y(N3390) );
  OR2X1 gate755 ( .A(N3007), .B(N2381), .Y(N3398) );
  OR2X1 gate756 ( .A(N3008), .B(N2382), .Y(N3404) );
  OR2X1 gate757 ( .A(N3009), .B(N2383), .Y(N3410) );
  OR2X1 gate758 ( .A(N3021), .B(N2397), .Y(N3416) );
  OR2X1 gate759 ( .A(N3022), .B(N2398), .Y(N3420) );
  OR2X1 gate760 ( .A(N3023), .B(N2399), .Y(N3424) );
  OR2X1 gate761 ( .A(N3024), .B(N2400), .Y(N3428) );
  OR2X1 gate762 ( .A(N3025), .B(N2401), .Y(N3432) );
  OR2X1 gate763 ( .A(N3026), .B(N2402), .Y(N3436) );
  OR2X1 gate764 ( .A(N3027), .B(N2403), .Y(N3440) );
  OR2X1 gate765 ( .A(N3028), .B(N2404), .Y(N3444) );
  OR2X1 gate766 ( .A(N3029), .B(N2405), .Y(N3448) );
  INVX1 gate767 ( .A(N2790), .Y(N3452) );
  INVX1 gate768 ( .A(N2793), .Y(N3453) );
  OR2X1 gate769 ( .A(N3034), .B(N2420), .Y(N3454) );
  OR2X1 gate770 ( .A(N3035), .B(N2421), .Y(N3458) );
  OR2X1 gate771 ( .A(N3036), .B(N2422), .Y(N3462) );
  OR2X1 gate772 ( .A(N3037), .B(N2423), .Y(N3466) );
  OR2X1 gate773 ( .A(N3038), .B(N2424), .Y(N3470) );
  OR2X1 gate774 ( .A(N3039), .B(N2425), .Y(N3474) );
  OR2X1 gate775 ( .A(N3040), .B(N2426), .Y(N3478) );
  OR2X1 gate776 ( .A(N3041), .B(N2427), .Y(N3482) );
  INVX1 gate777 ( .A(N2796), .Y(N3486) );
  BUFX2 gate778 ( .A(N2644), .Y(N3487) );
  BUFX2 gate779 ( .A(N2638), .Y(N3490) );
  BUFX2 gate780 ( .A(N2632), .Y(N3493) );
  BUFX2 gate781 ( .A(N2626), .Y(N3496) );
  BUFX2 gate782 ( .A(N2619), .Y(N3499) );
  BUFX2 gate783 ( .A(N2523), .Y(N3502) );
  NOR2X1 gate784 ( .A(N1167), .B(N2868), .Y(N3507) );
  BUFX2 gate785 ( .A(N2523), .Y(N3510) );
  NOR2X1 gate786 ( .A(N644), .B(N2619), .Y(N3515) );
  BUFX2 gate787 ( .A(N2644), .Y(N3518) );
  BUFX2 gate788 ( .A(N2638), .Y(N3521) );
  BUFX2 gate789 ( .A(N2632), .Y(N3524) );
  BUFX2 gate790 ( .A(N2626), .Y(N3527) );
  BUFX2 gate791 ( .A(N2619), .Y(N3530) );
  BUFX2 gate792 ( .A(N2619), .Y(N3535) );
  BUFX2 gate793 ( .A(N2632), .Y(N3539) );
  BUFX2 gate794 ( .A(N2626), .Y(N3542) );
  BUFX2 gate795 ( .A(N2644), .Y(N3545) );
  BUFX2 gate796 ( .A(N2638), .Y(N3548) );
  INVX1 gate797 ( .A(N2766), .Y(N3551) );
  INVX1 gate798 ( .A(N2769), .Y(N3552) );
  BUFX2 gate799 ( .A(N2442), .Y(N3553) );
  BUFX2 gate800 ( .A(N2450), .Y(N3557) );
  BUFX2 gate801 ( .A(N2446), .Y(N3560) );
  BUFX2 gate802 ( .A(N2458), .Y(N3563) );
  BUFX2 gate803 ( .A(N2454), .Y(N3566) );
  INVX1 gate804 ( .A(N2772), .Y(N3569) );
  INVX1 gate805 ( .A(N2775), .Y(N3570) );
  BUFX2 gate806 ( .A(N2554), .Y(N3571) );
  BUFX2 gate807 ( .A(N2567), .Y(N3574) );
  BUFX2 gate808 ( .A(N2561), .Y(N3577) );
  BUFX2 gate809 ( .A(N2482), .Y(N3580) );
  BUFX2 gate810 ( .A(N2573), .Y(N3583) );
  BUFX2 gate811 ( .A(N2496), .Y(N3586) );
  BUFX2 gate812 ( .A(N2488), .Y(N3589) );
  BUFX2 gate813 ( .A(N2508), .Y(N3592) );
  BUFX2 gate814 ( .A(N2502), .Y(N3595) );
  BUFX2 gate815 ( .A(N2508), .Y(N3598) );
  BUFX2 gate816 ( .A(N2502), .Y(N3601) );
  BUFX2 gate817 ( .A(N2496), .Y(N3604) );
  BUFX2 gate818 ( .A(N2482), .Y(N3607) );
  BUFX2 gate819 ( .A(N2573), .Y(N3610) );
  BUFX2 gate820 ( .A(N2567), .Y(N3613) );
  BUFX2 gate821 ( .A(N2561), .Y(N3616) );
  BUFX2 gate822 ( .A(N2488), .Y(N3619) );
  BUFX2 gate823 ( .A(N2554), .Y(N3622) );
  NOR2X1 gate824 ( .A(N734), .B(N2488), .Y(N3625) );
  NOR2X1 gate825 ( .A(N708), .B(N2554), .Y(N3628) );
  BUFX2 gate826 ( .A(N2508), .Y(N3631) );
  BUFX2 gate827 ( .A(N2502), .Y(N3634) );
  BUFX2 gate828 ( .A(N2496), .Y(N3637) );
  BUFX2 gate829 ( .A(N2488), .Y(N3640) );
  BUFX2 gate830 ( .A(N2482), .Y(N3643) );
  BUFX2 gate831 ( .A(N2573), .Y(N3646) );
  BUFX2 gate832 ( .A(N2567), .Y(N3649) );
  BUFX2 gate833 ( .A(N2561), .Y(N3652) );
  BUFX2 gate834 ( .A(N2554), .Y(N3655) );
  NOR2X1 gate835 ( .A(N2488), .B(N734), .Y(N3658) );
  BUFX2 gate836 ( .A(N2674), .Y(N3661) );
  BUFX2 gate837 ( .A(N2674), .Y(N3664) );
  BUFX2 gate838 ( .A(N2761), .Y(N3667) );
  BUFX2 gate839 ( .A(N2478), .Y(N3670) );
  BUFX2 gate840 ( .A(N2757), .Y(N3673) );
  BUFX2 gate841 ( .A(N2474), .Y(N3676) );
  BUFX2 gate842 ( .A(N2753), .Y(N3679) );
  BUFX2 gate843 ( .A(N2470), .Y(N3682) );
  BUFX2 gate844 ( .A(N2745), .Y(N3685) );
  BUFX2 gate845 ( .A(N2462), .Y(N3688) );
  BUFX2 gate846 ( .A(N2741), .Y(N3691) );
  BUFX2 gate847 ( .A(N2550), .Y(N3694) );
  BUFX2 gate848 ( .A(N2737), .Y(N3697) );
  BUFX2 gate849 ( .A(N2546), .Y(N3700) );
  BUFX2 gate850 ( .A(N2733), .Y(N3703) );
  BUFX2 gate851 ( .A(N2542), .Y(N3706) );
  BUFX2 gate852 ( .A(N2749), .Y(N3709) );
  BUFX2 gate853 ( .A(N2466), .Y(N3712) );
  BUFX2 gate854 ( .A(N2729), .Y(N3715) );
  BUFX2 gate855 ( .A(N2538), .Y(N3718) );
  BUFX2 gate856 ( .A(N2704), .Y(N3721) );
  BUFX2 gate857 ( .A(N2700), .Y(N3724) );
  BUFX2 gate858 ( .A(N2696), .Y(N3727) );
  BUFX2 gate859 ( .A(N2688), .Y(N3730) );
  BUFX2 gate860 ( .A(N2692), .Y(N3733) );
  BUFX2 gate861 ( .A(N2670), .Y(N3736) );
  BUFX2 gate862 ( .A(N2458), .Y(N3739) );
  BUFX2 gate863 ( .A(N2666), .Y(N3742) );
  BUFX2 gate864 ( .A(N2454), .Y(N3745) );
  BUFX2 gate865 ( .A(N2662), .Y(N3748) );
  BUFX2 gate866 ( .A(N2450), .Y(N3751) );
  BUFX2 gate867 ( .A(N2658), .Y(N3754) );
  BUFX2 gate868 ( .A(N2446), .Y(N3757) );
  BUFX2 gate869 ( .A(N2654), .Y(N3760) );
  BUFX2 gate870 ( .A(N2442), .Y(N3763) );
  BUFX2 gate871 ( .A(N2654), .Y(N3766) );
  BUFX2 gate872 ( .A(N2662), .Y(N3769) );
  BUFX2 gate873 ( .A(N2658), .Y(N3772) );
  BUFX2 gate874 ( .A(N2670), .Y(N3775) );
  BUFX2 gate875 ( .A(N2666), .Y(N3778) );
  INVX1 gate876 ( .A(N2784), .Y(N3781) );
  INVX1 gate877 ( .A(N2787), .Y(N3782) );
  OR2X1 gate878 ( .A(N2928), .B(N2326), .Y(N3783) );
  OR2X1 gate879 ( .A(N2933), .B(N2342), .Y(N3786) );
  OR2X1 gate880 ( .A(N2923), .B(N2321), .Y(N3789) );
  BUFX2 gate881 ( .A(N2688), .Y(N3792) );
  BUFX2 gate882 ( .A(N2696), .Y(N3795) );
  BUFX2 gate883 ( .A(N2692), .Y(N3798) );
  BUFX2 gate884 ( .A(N2704), .Y(N3801) );
  BUFX2 gate885 ( .A(N2700), .Y(N3804) );
  BUFX2 gate886 ( .A(N2604), .Y(N3807) );
  BUFX2 gate887 ( .A(N2611), .Y(N3810) );
  BUFX2 gate888 ( .A(N2607), .Y(N3813) );
  BUFX2 gate889 ( .A(N2615), .Y(N3816) );
  BUFX2 gate890 ( .A(N2538), .Y(N3819) );
  BUFX2 gate891 ( .A(N2546), .Y(N3822) );
  BUFX2 gate892 ( .A(N2542), .Y(N3825) );
  BUFX2 gate893 ( .A(N2462), .Y(N3828) );
  BUFX2 gate894 ( .A(N2550), .Y(N3831) );
  BUFX2 gate895 ( .A(N2470), .Y(N3834) );
  BUFX2 gate896 ( .A(N2466), .Y(N3837) );
  BUFX2 gate897 ( .A(N2478), .Y(N3840) );
  BUFX2 gate898 ( .A(N2474), .Y(N3843) );
  BUFX2 gate899 ( .A(N2615), .Y(N3846) );
  BUFX2 gate900 ( .A(N2611), .Y(N3849) );
  BUFX2 gate901 ( .A(N2607), .Y(N3852) );
  BUFX2 gate902 ( .A(N2680), .Y(N3855) );
  BUFX2 gate903 ( .A(N2729), .Y(N3858) );
  BUFX2 gate904 ( .A(N2737), .Y(N3861) );
  BUFX2 gate905 ( .A(N2733), .Y(N3864) );
  BUFX2 gate906 ( .A(N2745), .Y(N3867) );
  BUFX2 gate907 ( .A(N2741), .Y(N3870) );
  BUFX2 gate908 ( .A(N2753), .Y(N3873) );
  BUFX2 gate909 ( .A(N2749), .Y(N3876) );
  BUFX2 gate910 ( .A(N2761), .Y(N3879) );
  BUFX2 gate911 ( .A(N2757), .Y(N3882) );
  OR2X1 gate912 ( .A(N3033), .B(N2419), .Y(N3885) );
  OR2X1 gate913 ( .A(N3032), .B(N2418), .Y(N3888) );
  OR2X1 gate914 ( .A(N3020), .B(N2396), .Y(N3891) );
  NAND2X1 gate915 ( .A(N3067), .B(N2117), .Y(N3953) );
  INVX1 gate916 ( .A(N3067), .Y(N3954) );
  NAND2X1 gate917 ( .A(N3070), .B(N2537), .Y(N3955) );
  INVX1 gate918 ( .A(N3070), .Y(N3956) );
  INVX1 gate919 ( .A(N3073), .Y(N3958) );
  INVX1 gate920 ( .A(N3080), .Y(N3964) );
  OR2X1 gate921 ( .A(N1649), .B(N3379), .Y(N4193) );
  OR2X1 gate922_1 ( .A(N1167), .B(N2867), .Y(N4303_1) );
  OR2X1 gate922 ( .A(N3130), .B(N4303_1), .Y(N4303) );
  INVX1 gate923 ( .A(N3061), .Y(N4308) );
  INVX1 gate924 ( .A(N3064), .Y(N4313) );
  NAND2X1 gate925 ( .A(N2769), .B(N3551), .Y(N4326) );
  NAND2X1 gate926 ( .A(N2766), .B(N3552), .Y(N4327) );
  NAND2X1 gate927 ( .A(N2775), .B(N3569), .Y(N4333) );
  NAND2X1 gate928 ( .A(N2772), .B(N3570), .Y(N4334) );
  NAND2X1 gate929 ( .A(N2787), .B(N3781), .Y(N4411) );
  NAND2X1 gate930 ( .A(N2784), .B(N3782), .Y(N4412) );
  NAND2X1 gate931 ( .A(N3487), .B(N1828), .Y(N4463) );
  INVX1 gate932 ( .A(N3487), .Y(N4464) );
  NAND2X1 gate933 ( .A(N3490), .B(N1829), .Y(N4465) );
  INVX1 gate934 ( .A(N3490), .Y(N4466) );
  NAND2X1 gate935 ( .A(N3493), .B(N2267), .Y(N4467) );
  INVX1 gate936 ( .A(N3493), .Y(N4468) );
  NAND2X1 gate937 ( .A(N3496), .B(N1830), .Y(N4469) );
  INVX1 gate938 ( .A(N3496), .Y(N4470) );
  NAND2X1 gate939 ( .A(N3499), .B(N1833), .Y(N4471) );
  INVX1 gate940 ( .A(N3499), .Y(N4472) );
  INVX1 gate941 ( .A(N3122), .Y(N4473) );
  INVX1 gate942 ( .A(N3126), .Y(N4474) );
  NAND2X1 gate943 ( .A(N3518), .B(N1840), .Y(N4475) );
  INVX1 gate944 ( .A(N3518), .Y(N4476) );
  NAND2X1 gate945 ( .A(N3521), .B(N1841), .Y(N4477) );
  INVX1 gate946 ( .A(N3521), .Y(N4478) );
  NAND2X1 gate947 ( .A(N3524), .B(N2275), .Y(N4479) );
  INVX1 gate948 ( .A(N3524), .Y(N4480) );
  NAND2X1 gate949 ( .A(N3527), .B(N1842), .Y(N4481) );
  INVX1 gate950 ( .A(N3527), .Y(N4482) );
  NAND2X1 gate951 ( .A(N3530), .B(N1843), .Y(N4483) );
  INVX1 gate952 ( .A(N3530), .Y(N4484) );
  INVX1 gate953 ( .A(N3155), .Y(N4485) );
  INVX1 gate954 ( .A(N3159), .Y(N4486) );
  NAND2X1 gate955 ( .A(N1721), .B(N3954), .Y(N4487) );
  NAND2X1 gate956 ( .A(N2235), .B(N3956), .Y(N4488) );
  INVX1 gate957 ( .A(N3535), .Y(N4489) );
  NAND2X1 gate958 ( .A(N3535), .B(N3958), .Y(N4490) );
  INVX1 gate959 ( .A(N3539), .Y(N4491) );
  INVX1 gate960 ( .A(N3542), .Y(N4492) );
  INVX1 gate961 ( .A(N3545), .Y(N4493) );
  INVX1 gate962 ( .A(N3548), .Y(N4494) );
  INVX1 gate963 ( .A(N3553), .Y(N4495) );
  NAND2X1 gate964 ( .A(N3553), .B(N3964), .Y(N4496) );
  INVX1 gate965 ( .A(N3557), .Y(N4497) );
  INVX1 gate966 ( .A(N3560), .Y(N4498) );
  INVX1 gate967 ( .A(N3563), .Y(N4499) );
  INVX1 gate968 ( .A(N3566), .Y(N4500) );
  INVX1 gate969 ( .A(N3571), .Y(N4501) );
  NAND2X1 gate970 ( .A(N3571), .B(N3167), .Y(N4502) );
  INVX1 gate971 ( .A(N3574), .Y(N4503) );
  INVX1 gate972 ( .A(N3577), .Y(N4504) );
  INVX1 gate973 ( .A(N3580), .Y(N4505) );
  INVX1 gate974 ( .A(N3583), .Y(N4506) );
  NAND2X1 gate975 ( .A(N3598), .B(N1867), .Y(N4507) );
  INVX1 gate976 ( .A(N3598), .Y(N4508) );
  NAND2X1 gate977 ( .A(N3601), .B(N1868), .Y(N4509) );
  INVX1 gate978 ( .A(N3601), .Y(N4510) );
  NAND2X1 gate979 ( .A(N3604), .B(N1869), .Y(N4511) );
  INVX1 gate980 ( .A(N3604), .Y(N4512) );
  NAND2X1 gate981 ( .A(N3607), .B(N1870), .Y(N4513) );
  INVX1 gate982 ( .A(N3607), .Y(N4514) );
  NAND2X1 gate983 ( .A(N3610), .B(N1871), .Y(N4515) );
  INVX1 gate984 ( .A(N3610), .Y(N4516) );
  NAND2X1 gate985 ( .A(N3613), .B(N1872), .Y(N4517) );
  INVX1 gate986 ( .A(N3613), .Y(N4518) );
  NAND2X1 gate987 ( .A(N3616), .B(N1873), .Y(N4519) );
  INVX1 gate988 ( .A(N3616), .Y(N4520) );
  NAND2X1 gate989 ( .A(N3619), .B(N1874), .Y(N4521) );
  INVX1 gate990 ( .A(N3619), .Y(N4522) );
  NAND2X1 gate991 ( .A(N3622), .B(N1875), .Y(N4523) );
  INVX1 gate992 ( .A(N3622), .Y(N4524) );
  NAND2X1 gate993 ( .A(N3631), .B(N1876), .Y(N4525) );
  INVX1 gate994 ( .A(N3631), .Y(N4526) );
  NAND2X1 gate995 ( .A(N3634), .B(N1877), .Y(N4527) );
  INVX1 gate996 ( .A(N3634), .Y(N4528) );
  NAND2X1 gate997 ( .A(N3637), .B(N1878), .Y(N4529) );
  INVX1 gate998 ( .A(N3637), .Y(N4530) );
  NAND2X1 gate999 ( .A(N3640), .B(N1879), .Y(N4531) );
  INVX1 gate1000 ( .A(N3640), .Y(N4532) );
  NAND2X1 gate1001 ( .A(N3643), .B(N1880), .Y(N4533) );
  INVX1 gate1002 ( .A(N3643), .Y(N4534) );
  NAND2X1 gate1003 ( .A(N3646), .B(N1881), .Y(N4535) );
  INVX1 gate1004 ( .A(N3646), .Y(N4536) );
  NAND2X1 gate1005 ( .A(N3649), .B(N1882), .Y(N4537) );
  INVX1 gate1006 ( .A(N3649), .Y(N4538) );
  NAND2X1 gate1007 ( .A(N3652), .B(N1883), .Y(N4539) );
  INVX1 gate1008 ( .A(N3652), .Y(N4540) );
  NAND2X1 gate1009 ( .A(N3655), .B(N1884), .Y(N4541) );
  INVX1 gate1010 ( .A(N3655), .Y(N4542) );
  INVX1 gate1011 ( .A(N3658), .Y(N4543) );
  AND2X1 gate1012 ( .A(N806), .B(N3293), .Y(N4544) );
  AND2X1 gate1013 ( .A(N800), .B(N3287), .Y(N4545) );
  AND2X1 gate1014 ( .A(N794), .B(N3281), .Y(N4549) );
  AND2X1 gate1015 ( .A(N3273), .B(N786), .Y(N4555) );
  AND2X1 gate1016 ( .A(N780), .B(N3267), .Y(N4562) );
  AND2X1 gate1017 ( .A(N774), .B(N3355), .Y(N4563) );
  AND2X1 gate1018 ( .A(N768), .B(N3349), .Y(N4566) );
  AND2X1 gate1019 ( .A(N762), .B(N3343), .Y(N4570) );
  INVX1 gate1020 ( .A(N3661), .Y(N4575) );
  AND2X1 gate1021 ( .A(N806), .B(N3293), .Y(N4576) );
  AND2X1 gate1022 ( .A(N800), .B(N3287), .Y(N4577) );
  AND2X1 gate1023 ( .A(N794), .B(N3281), .Y(N4581) );
  AND2X1 gate1024 ( .A(N786), .B(N3273), .Y(N4586) );
  AND2X1 gate1025 ( .A(N780), .B(N3267), .Y(N4592) );
  AND2X1 gate1026 ( .A(N774), .B(N3355), .Y(N4593) );
  AND2X1 gate1027 ( .A(N768), .B(N3349), .Y(N4597) );
  AND2X1 gate1028 ( .A(N762), .B(N3343), .Y(N4603) );
  INVX1 gate1029 ( .A(N3664), .Y(N4610) );
  INVX1 gate1030 ( .A(N3667), .Y(N4611) );
  INVX1 gate1031 ( .A(N3670), .Y(N4612) );
  INVX1 gate1032 ( .A(N3673), .Y(N4613) );
  INVX1 gate1033 ( .A(N3676), .Y(N4614) );
  INVX1 gate1034 ( .A(N3679), .Y(N4615) );
  INVX1 gate1035 ( .A(N3682), .Y(N4616) );
  INVX1 gate1036 ( .A(N3685), .Y(N4617) );
  INVX1 gate1037 ( .A(N3688), .Y(N4618) );
  INVX1 gate1038 ( .A(N3691), .Y(N4619) );
  INVX1 gate1039 ( .A(N3694), .Y(N4620) );
  INVX1 gate1040 ( .A(N3697), .Y(N4621) );
  INVX1 gate1041 ( .A(N3700), .Y(N4622) );
  INVX1 gate1042 ( .A(N3703), .Y(N4623) );
  INVX1 gate1043 ( .A(N3706), .Y(N4624) );
  INVX1 gate1044 ( .A(N3709), .Y(N4625) );
  INVX1 gate1045 ( .A(N3712), .Y(N4626) );
  INVX1 gate1046 ( .A(N3715), .Y(N4627) );
  INVX1 gate1047 ( .A(N3718), .Y(N4628) );
  INVX1 gate1048 ( .A(N3721), .Y(N4629) );
  AND2X1 gate1049 ( .A(N3448), .B(N2704), .Y(N4630) );
  INVX1 gate1050 ( .A(N3724), .Y(N4631) );
  AND2X1 gate1051 ( .A(N3444), .B(N2700), .Y(N4632) );
  INVX1 gate1052 ( .A(N3727), .Y(N4633) );
  AND2X1 gate1053 ( .A(N3440), .B(N2696), .Y(N4634) );
  AND2X1 gate1054 ( .A(N3436), .B(N2692), .Y(N4635) );
  INVX1 gate1055 ( .A(N3730), .Y(N4636) );
  AND2X1 gate1056 ( .A(N3432), .B(N2688), .Y(N4637) );
  AND2X1 gate1057 ( .A(N3428), .B(N3311), .Y(N4638) );
  AND2X1 gate1058 ( .A(N3424), .B(N3307), .Y(N4639) );
  AND2X1 gate1059 ( .A(N3420), .B(N3303), .Y(N4640) );
  AND2X1 gate1060 ( .A(N3416), .B(N3299), .Y(N4641) );
  INVX1 gate1061 ( .A(N3733), .Y(N4642) );
  INVX1 gate1062 ( .A(N3736), .Y(N4643) );
  INVX1 gate1063 ( .A(N3739), .Y(N4644) );
  INVX1 gate1064 ( .A(N3742), .Y(N4645) );
  INVX1 gate1065 ( .A(N3745), .Y(N4646) );
  INVX1 gate1066 ( .A(N3748), .Y(N4647) );
  INVX1 gate1067 ( .A(N3751), .Y(N4648) );
  INVX1 gate1068 ( .A(N3754), .Y(N4649) );
  INVX1 gate1069 ( .A(N3757), .Y(N4650) );
  INVX1 gate1070 ( .A(N3760), .Y(N4651) );
  INVX1 gate1071 ( .A(N3763), .Y(N4652) );
  INVX1 gate1072 ( .A(N3375), .Y(N4653) );
  AND2X1 gate1073 ( .A(N865), .B(N3410), .Y(N4656) );
  AND2X1 gate1074 ( .A(N859), .B(N3404), .Y(N4657) );
  AND2X1 gate1075 ( .A(N853), .B(N3398), .Y(N4661) );
  AND2X1 gate1076 ( .A(N3390), .B(N845), .Y(N4667) );
  AND2X1 gate1077 ( .A(N839), .B(N3384), .Y(N4674) );
  AND2X1 gate1078 ( .A(N833), .B(N3334), .Y(N4675) );
  AND2X1 gate1079 ( .A(N827), .B(N3328), .Y(N4678) );
  AND2X1 gate1080 ( .A(N821), .B(N3322), .Y(N4682) );
  AND2X1 gate1081 ( .A(N814), .B(N3315), .Y(N4687) );
  INVX1 gate1082 ( .A(N3766), .Y(N4693) );
  NAND2X1 gate1083 ( .A(N3766), .B(N3380), .Y(N4694) );
  INVX1 gate1084 ( .A(N3769), .Y(N4695) );
  INVX1 gate1085 ( .A(N3772), .Y(N4696) );
  INVX1 gate1086 ( .A(N3775), .Y(N4697) );
  INVX1 gate1087 ( .A(N3778), .Y(N4698) );
  INVX1 gate1088 ( .A(N3783), .Y(N4699) );
  INVX1 gate1089 ( .A(N3786), .Y(N4700) );
  AND2X1 gate1090 ( .A(N865), .B(N3410), .Y(N4701) );
  AND2X1 gate1091 ( .A(N859), .B(N3404), .Y(N4702) );
  AND2X1 gate1092 ( .A(N853), .B(N3398), .Y(N4706) );
  AND2X1 gate1093 ( .A(N845), .B(N3390), .Y(N4711) );
  AND2X1 gate1094 ( .A(N839), .B(N3384), .Y(N4717) );
  AND2X1 gate1095 ( .A(N833), .B(N3334), .Y(N4718) );
  AND2X1 gate1096 ( .A(N827), .B(N3328), .Y(N4722) );
  AND2X1 gate1097 ( .A(N821), .B(N3322), .Y(N4728) );
  AND2X1 gate1098 ( .A(N814), .B(N3315), .Y(N4735) );
  INVX1 gate1099 ( .A(N3789), .Y(N4743) );
  INVX1 gate1100 ( .A(N3792), .Y(N4744) );
  INVX1 gate1101 ( .A(N3807), .Y(N4745) );
  NAND2X1 gate1102 ( .A(N3807), .B(N3452), .Y(N4746) );
  INVX1 gate1103 ( .A(N3810), .Y(N4747) );
  INVX1 gate1104 ( .A(N3813), .Y(N4748) );
  INVX1 gate1105 ( .A(N3816), .Y(N4749) );
  INVX1 gate1106 ( .A(N3819), .Y(N4750) );
  NAND2X1 gate1107 ( .A(N3819), .B(N3453), .Y(N4751) );
  INVX1 gate1108 ( .A(N3822), .Y(N4752) );
  INVX1 gate1109 ( .A(N3825), .Y(N4753) );
  INVX1 gate1110 ( .A(N3828), .Y(N4754) );
  INVX1 gate1111 ( .A(N3831), .Y(N4755) );
  AND2X1 gate1112 ( .A(N3482), .B(N3263), .Y(N4756) );
  AND2X1 gate1113 ( .A(N3478), .B(N3259), .Y(N4757) );
  AND2X1 gate1114 ( .A(N3474), .B(N3255), .Y(N4758) );
  AND2X1 gate1115 ( .A(N3470), .B(N3251), .Y(N4759) );
  AND2X1 gate1116 ( .A(N3466), .B(N3247), .Y(N4760) );
  INVX1 gate1117 ( .A(N3846), .Y(N4761) );
  AND2X1 gate1118 ( .A(N3462), .B(N2615), .Y(N4762) );
  INVX1 gate1119 ( .A(N3849), .Y(N4763) );
  AND2X1 gate1120 ( .A(N3458), .B(N2611), .Y(N4764) );
  INVX1 gate1121 ( .A(N3852), .Y(N4765) );
  AND2X1 gate1122 ( .A(N3454), .B(N2607), .Y(N4766) );
  AND2X1 gate1123 ( .A(N2680), .B(N3381), .Y(N4767) );
  INVX1 gate1124 ( .A(N3855), .Y(N4768) );
  AND2X1 gate1125 ( .A(N3340), .B(N695), .Y(N4769) );
  INVX1 gate1126 ( .A(N3858), .Y(N4775) );
  NAND2X1 gate1127 ( .A(N3858), .B(N3486), .Y(N4776) );
  INVX1 gate1128 ( .A(N3861), .Y(N4777) );
  INVX1 gate1129 ( .A(N3864), .Y(N4778) );
  INVX1 gate1130 ( .A(N3867), .Y(N4779) );
  INVX1 gate1131 ( .A(N3870), .Y(N4780) );
  INVX1 gate1132 ( .A(N3885), .Y(N4781) );
  INVX1 gate1133 ( .A(N3888), .Y(N4782) );
  INVX1 gate1134 ( .A(N3891), .Y(N4783) );
  OR2X1 gate1135 ( .A(N3131), .B(N3134), .Y(N4784) );
  INVX1 gate1136 ( .A(N3502), .Y(N4789) );
  INVX1 gate1137 ( .A(N3131), .Y(N4790) );
  INVX1 gate1138 ( .A(N3507), .Y(N4793) );
  INVX1 gate1139 ( .A(N3510), .Y(N4794) );
  INVX1 gate1140 ( .A(N3515), .Y(N4795) );
  BUFX2 gate1141 ( .A(N3114), .Y(N4796) );
  INVX1 gate1142 ( .A(N3586), .Y(N4799) );
  INVX1 gate1143 ( .A(N3589), .Y(N4800) );
  INVX1 gate1144 ( .A(N3592), .Y(N4801) );
  INVX1 gate1145 ( .A(N3595), .Y(N4802) );
  NAND2X1 gate1146 ( .A(N4326), .B(N4327), .Y(N4803) );
  NAND2X1 gate1147 ( .A(N4333), .B(N4334), .Y(N4806) );
  INVX1 gate1148 ( .A(N3625), .Y(N4809) );
  BUFX2 gate1149 ( .A(N3178), .Y(N4810) );
  INVX1 gate1150 ( .A(N3628), .Y(N4813) );
  BUFX2 gate1151 ( .A(N3202), .Y(N4814) );
  BUFX2 gate1152 ( .A(N3221), .Y(N4817) );
  BUFX2 gate1153 ( .A(N3293), .Y(N4820) );
  BUFX2 gate1154 ( .A(N3287), .Y(N4823) );
  BUFX2 gate1155 ( .A(N3281), .Y(N4826) );
  BUFX2 gate1156 ( .A(N3273), .Y(N4829) );
  BUFX2 gate1157 ( .A(N3267), .Y(N4832) );
  BUFX2 gate1158 ( .A(N3355), .Y(N4835) );
  BUFX2 gate1159 ( .A(N3349), .Y(N4838) );
  BUFX2 gate1160 ( .A(N3343), .Y(N4841) );
  NOR2X1 gate1161 ( .A(N3273), .B(N786), .Y(N4844) );
  BUFX2 gate1162 ( .A(N3293), .Y(N4847) );
  BUFX2 gate1163 ( .A(N3287), .Y(N4850) );
  BUFX2 gate1164 ( .A(N3281), .Y(N4853) );
  BUFX2 gate1165 ( .A(N3267), .Y(N4856) );
  BUFX2 gate1166 ( .A(N3355), .Y(N4859) );
  BUFX2 gate1167 ( .A(N3349), .Y(N4862) );
  BUFX2 gate1168 ( .A(N3343), .Y(N4865) );
  BUFX2 gate1169 ( .A(N3273), .Y(N4868) );
  NOR2X1 gate1170 ( .A(N786), .B(N3273), .Y(N4871) );
  BUFX2 gate1171 ( .A(N3448), .Y(N4874) );
  BUFX2 gate1172 ( .A(N3444), .Y(N4877) );
  BUFX2 gate1173 ( .A(N3440), .Y(N4880) );
  BUFX2 gate1174 ( .A(N3432), .Y(N4883) );
  BUFX2 gate1175 ( .A(N3428), .Y(N4886) );
  BUFX2 gate1176 ( .A(N3311), .Y(N4889) );
  BUFX2 gate1177 ( .A(N3424), .Y(N4892) );
  BUFX2 gate1178 ( .A(N3307), .Y(N4895) );
  BUFX2 gate1179 ( .A(N3420), .Y(N4898) );
  BUFX2 gate1180 ( .A(N3303), .Y(N4901) );
  BUFX2 gate1181 ( .A(N3436), .Y(N4904) );
  BUFX2 gate1182 ( .A(N3416), .Y(N4907) );
  BUFX2 gate1183 ( .A(N3299), .Y(N4910) );
  BUFX2 gate1184 ( .A(N3410), .Y(N4913) );
  BUFX2 gate1185 ( .A(N3404), .Y(N4916) );
  BUFX2 gate1186 ( .A(N3398), .Y(N4919) );
  BUFX2 gate1187 ( .A(N3390), .Y(N4922) );
  BUFX2 gate1188 ( .A(N3384), .Y(N4925) );
  BUFX2 gate1189 ( .A(N3334), .Y(N4928) );
  BUFX2 gate1190 ( .A(N3328), .Y(N4931) );
  BUFX2 gate1191 ( .A(N3322), .Y(N4934) );
  BUFX2 gate1192 ( .A(N3315), .Y(N4937) );
  NOR2X1 gate1193 ( .A(N3390), .B(N845), .Y(N4940) );
  BUFX2 gate1194 ( .A(N3315), .Y(N4943) );
  BUFX2 gate1195 ( .A(N3328), .Y(N4946) );
  BUFX2 gate1196 ( .A(N3322), .Y(N4949) );
  BUFX2 gate1197 ( .A(N3384), .Y(N4952) );
  BUFX2 gate1198 ( .A(N3334), .Y(N4955) );
  BUFX2 gate1199 ( .A(N3398), .Y(N4958) );
  BUFX2 gate1200 ( .A(N3390), .Y(N4961) );
  BUFX2 gate1201 ( .A(N3410), .Y(N4964) );
  BUFX2 gate1202 ( .A(N3404), .Y(N4967) );
  BUFX2 gate1203 ( .A(N3340), .Y(N4970) );
  BUFX2 gate1204 ( .A(N3349), .Y(N4973) );
  BUFX2 gate1205 ( .A(N3343), .Y(N4976) );
  BUFX2 gate1206 ( .A(N3267), .Y(N4979) );
  BUFX2 gate1207 ( .A(N3355), .Y(N4982) );
  BUFX2 gate1208 ( .A(N3281), .Y(N4985) );
  BUFX2 gate1209 ( .A(N3273), .Y(N4988) );
  BUFX2 gate1210 ( .A(N3293), .Y(N4991) );
  BUFX2 gate1211 ( .A(N3287), .Y(N4994) );
  NAND2X1 gate1212 ( .A(N4411), .B(N4412), .Y(N4997) );
  BUFX2 gate1213 ( .A(N3410), .Y(N5000) );
  BUFX2 gate1214 ( .A(N3404), .Y(N5003) );
  BUFX2 gate1215 ( .A(N3398), .Y(N5006) );
  BUFX2 gate1216 ( .A(N3384), .Y(N5009) );
  BUFX2 gate1217 ( .A(N3334), .Y(N5012) );
  BUFX2 gate1218 ( .A(N3328), .Y(N5015) );
  BUFX2 gate1219 ( .A(N3322), .Y(N5018) );
  BUFX2 gate1220 ( .A(N3390), .Y(N5021) );
  BUFX2 gate1221 ( .A(N3315), .Y(N5024) );
  NOR2X1 gate1222 ( .A(N845), .B(N3390), .Y(N5027) );
  NOR2X1 gate1223 ( .A(N814), .B(N3315), .Y(N5030) );
  BUFX2 gate1224 ( .A(N3299), .Y(N5033) );
  BUFX2 gate1225 ( .A(N3307), .Y(N5036) );
  BUFX2 gate1226 ( .A(N3303), .Y(N5039) );
  BUFX2 gate1227 ( .A(N3311), .Y(N5042) );
  INVX1 gate1228 ( .A(N3795), .Y(N5045) );
  INVX1 gate1229 ( .A(N3798), .Y(N5046) );
  INVX1 gate1230 ( .A(N3801), .Y(N5047) );
  INVX1 gate1231 ( .A(N3804), .Y(N5048) );
  BUFX2 gate1232 ( .A(N3247), .Y(N5049) );
  BUFX2 gate1233 ( .A(N3255), .Y(N5052) );
  BUFX2 gate1234 ( .A(N3251), .Y(N5055) );
  BUFX2 gate1235 ( .A(N3263), .Y(N5058) );
  BUFX2 gate1236 ( .A(N3259), .Y(N5061) );
  INVX1 gate1237 ( .A(N3834), .Y(N5064) );
  INVX1 gate1238 ( .A(N3837), .Y(N5065) );
  INVX1 gate1239 ( .A(N3840), .Y(N5066) );
  INVX1 gate1240 ( .A(N3843), .Y(N5067) );
  BUFX2 gate1241 ( .A(N3482), .Y(N5068) );
  BUFX2 gate1242 ( .A(N3263), .Y(N5071) );
  BUFX2 gate1243 ( .A(N3478), .Y(N5074) );
  BUFX2 gate1244 ( .A(N3259), .Y(N5077) );
  BUFX2 gate1245 ( .A(N3474), .Y(N5080) );
  BUFX2 gate1246 ( .A(N3255), .Y(N5083) );
  BUFX2 gate1247 ( .A(N3466), .Y(N5086) );
  BUFX2 gate1248 ( .A(N3247), .Y(N5089) );
  BUFX2 gate1249 ( .A(N3462), .Y(N5092) );
  BUFX2 gate1250 ( .A(N3458), .Y(N5095) );
  BUFX2 gate1251 ( .A(N3454), .Y(N5098) );
  BUFX2 gate1252 ( .A(N3470), .Y(N5101) );
  BUFX2 gate1253 ( .A(N3251), .Y(N5104) );
  BUFX2 gate1254 ( .A(N3381), .Y(N5107) );
  INVX1 gate1255 ( .A(N3873), .Y(N5110) );
  INVX1 gate1256 ( .A(N3876), .Y(N5111) );
  INVX1 gate1257 ( .A(N3879), .Y(N5112) );
  INVX1 gate1258 ( .A(N3882), .Y(N5113) );
  BUFX2 gate1259 ( .A(N3458), .Y(N5114) );
  BUFX2 gate1260 ( .A(N3454), .Y(N5117) );
  BUFX2 gate1261 ( .A(N3466), .Y(N5120) );
  BUFX2 gate1262 ( .A(N3462), .Y(N5123) );
  BUFX2 gate1263 ( .A(N3474), .Y(N5126) );
  BUFX2 gate1264 ( .A(N3470), .Y(N5129) );
  BUFX2 gate1265 ( .A(N3482), .Y(N5132) );
  BUFX2 gate1266 ( .A(N3478), .Y(N5135) );
  BUFX2 gate1267 ( .A(N3416), .Y(N5138) );
  BUFX2 gate1268 ( .A(N3424), .Y(N5141) );
  BUFX2 gate1269 ( .A(N3420), .Y(N5144) );
  BUFX2 gate1270 ( .A(N3432), .Y(N5147) );
  BUFX2 gate1271 ( .A(N3428), .Y(N5150) );
  BUFX2 gate1272 ( .A(N3440), .Y(N5153) );
  BUFX2 gate1273 ( .A(N3436), .Y(N5156) );
  BUFX2 gate1274 ( .A(N3448), .Y(N5159) );
  BUFX2 gate1275 ( .A(N3444), .Y(N5162) );
  NAND2X1 gate1276 ( .A(N4486), .B(N4485), .Y(N5165) );
  NAND2X1 gate1277 ( .A(N4474), .B(N4473), .Y(N5166) );
  NAND2X1 gate1278 ( .A(N1290), .B(N4464), .Y(N5167) );
  NAND2X1 gate1279 ( .A(N1293), .B(N4466), .Y(N5168) );
  NAND2X1 gate1280 ( .A(N2074), .B(N4468), .Y(N5169) );
  NAND2X1 gate1281 ( .A(N1296), .B(N4470), .Y(N5170) );
  NAND2X1 gate1282 ( .A(N1302), .B(N4472), .Y(N5171) );
  NAND2X1 gate1283 ( .A(N1314), .B(N4476), .Y(N5172) );
  NAND2X1 gate1284 ( .A(N1317), .B(N4478), .Y(N5173) );
  NAND2X1 gate1285 ( .A(N2081), .B(N4480), .Y(N5174) );
  NAND2X1 gate1286 ( .A(N1320), .B(N4482), .Y(N5175) );
  NAND2X1 gate1287 ( .A(N1323), .B(N4484), .Y(N5176) );
  NAND2X1 gate1288 ( .A(N3953), .B(N4487), .Y(N5177) );
  NAND2X1 gate1289 ( .A(N3955), .B(N4488), .Y(N5178) );
  NAND2X1 gate1290 ( .A(N3073), .B(N4489), .Y(N5179) );
  NAND2X1 gate1291 ( .A(N3542), .B(N4491), .Y(N5180) );
  NAND2X1 gate1292 ( .A(N3539), .B(N4492), .Y(N5181) );
  NAND2X1 gate1293 ( .A(N3548), .B(N4493), .Y(N5182) );
  NAND2X1 gate1294 ( .A(N3545), .B(N4494), .Y(N5183) );
  NAND2X1 gate1295 ( .A(N3080), .B(N4495), .Y(N5184) );
  NAND2X1 gate1296 ( .A(N3560), .B(N4497), .Y(N5185) );
  NAND2X1 gate1297 ( .A(N3557), .B(N4498), .Y(N5186) );
  NAND2X1 gate1298 ( .A(N3566), .B(N4499), .Y(N5187) );
  NAND2X1 gate1299 ( .A(N3563), .B(N4500), .Y(N5188) );
  NAND2X1 gate1300 ( .A(N2778), .B(N4501), .Y(N5189) );
  NAND2X1 gate1301 ( .A(N3577), .B(N4503), .Y(N5190) );
  NAND2X1 gate1302 ( .A(N3574), .B(N4504), .Y(N5191) );
  NAND2X1 gate1303 ( .A(N3583), .B(N4505), .Y(N5192) );
  NAND2X1 gate1304 ( .A(N3580), .B(N4506), .Y(N5193) );
  NAND2X1 gate1305 ( .A(N1326), .B(N4508), .Y(N5196) );
  NAND2X1 gate1306 ( .A(N1329), .B(N4510), .Y(N5197) );
  NAND2X1 gate1307 ( .A(N1332), .B(N4512), .Y(N5198) );
  NAND2X1 gate1308 ( .A(N1335), .B(N4514), .Y(N5199) );
  NAND2X1 gate1309 ( .A(N1338), .B(N4516), .Y(N5200) );
  NAND2X1 gate1310 ( .A(N1341), .B(N4518), .Y(N5201) );
  NAND2X1 gate1311 ( .A(N1344), .B(N4520), .Y(N5202) );
  NAND2X1 gate1312 ( .A(N1347), .B(N4522), .Y(N5203) );
  NAND2X1 gate1313 ( .A(N1350), .B(N4524), .Y(N5204) );
  NAND2X1 gate1314 ( .A(N1353), .B(N4526), .Y(N5205) );
  NAND2X1 gate1315 ( .A(N1356), .B(N4528), .Y(N5206) );
  NAND2X1 gate1316 ( .A(N1359), .B(N4530), .Y(N5207) );
  NAND2X1 gate1317 ( .A(N1362), .B(N4532), .Y(N5208) );
  NAND2X1 gate1318 ( .A(N1365), .B(N4534), .Y(N5209) );
  NAND2X1 gate1319 ( .A(N1368), .B(N4536), .Y(N5210) );
  NAND2X1 gate1320 ( .A(N1371), .B(N4538), .Y(N5211) );
  NAND2X1 gate1321 ( .A(N1374), .B(N4540), .Y(N5212) );
  NAND2X1 gate1322 ( .A(N1377), .B(N4542), .Y(N5213) );
  NAND2X1 gate1323 ( .A(N3670), .B(N4611), .Y(N5283) );
  NAND2X1 gate1324 ( .A(N3667), .B(N4612), .Y(N5284) );
  NAND2X1 gate1325 ( .A(N3676), .B(N4613), .Y(N5285) );
  NAND2X1 gate1326 ( .A(N3673), .B(N4614), .Y(N5286) );
  NAND2X1 gate1327 ( .A(N3682), .B(N4615), .Y(N5287) );
  NAND2X1 gate1328 ( .A(N3679), .B(N4616), .Y(N5288) );
  NAND2X1 gate1329 ( .A(N3688), .B(N4617), .Y(N5289) );
  NAND2X1 gate1330 ( .A(N3685), .B(N4618), .Y(N5290) );
  NAND2X1 gate1331 ( .A(N3694), .B(N4619), .Y(N5291) );
  NAND2X1 gate1332 ( .A(N3691), .B(N4620), .Y(N5292) );
  NAND2X1 gate1333 ( .A(N3700), .B(N4621), .Y(N5293) );
  NAND2X1 gate1334 ( .A(N3697), .B(N4622), .Y(N5294) );
  NAND2X1 gate1335 ( .A(N3706), .B(N4623), .Y(N5295) );
  NAND2X1 gate1336 ( .A(N3703), .B(N4624), .Y(N5296) );
  NAND2X1 gate1337 ( .A(N3712), .B(N4625), .Y(N5297) );
  NAND2X1 gate1338 ( .A(N3709), .B(N4626), .Y(N5298) );
  NAND2X1 gate1339 ( .A(N3718), .B(N4627), .Y(N5299) );
  NAND2X1 gate1340 ( .A(N3715), .B(N4628), .Y(N5300) );
  NAND2X1 gate1341 ( .A(N3739), .B(N4643), .Y(N5314) );
  NAND2X1 gate1342 ( .A(N3736), .B(N4644), .Y(N5315) );
  NAND2X1 gate1343 ( .A(N3745), .B(N4645), .Y(N5316) );
  NAND2X1 gate1344 ( .A(N3742), .B(N4646), .Y(N5317) );
  NAND2X1 gate1345 ( .A(N3751), .B(N4647), .Y(N5318) );
  NAND2X1 gate1346 ( .A(N3748), .B(N4648), .Y(N5319) );
  NAND2X1 gate1347 ( .A(N3757), .B(N4649), .Y(N5320) );
  NAND2X1 gate1348 ( .A(N3754), .B(N4650), .Y(N5321) );
  NAND2X1 gate1349 ( .A(N3763), .B(N4651), .Y(N5322) );
  NAND2X1 gate1350 ( .A(N3760), .B(N4652), .Y(N5323) );
  INVX1 gate1351 ( .A(N4193), .Y(N5324) );
  NAND2X1 gate1352 ( .A(N2781), .B(N4693), .Y(N5363) );
  NAND2X1 gate1353 ( .A(N3772), .B(N4695), .Y(N5364) );
  NAND2X1 gate1354 ( .A(N3769), .B(N4696), .Y(N5365) );
  NAND2X1 gate1355 ( .A(N3778), .B(N4697), .Y(N5366) );
  NAND2X1 gate1356 ( .A(N3775), .B(N4698), .Y(N5367) );
  NAND2X1 gate1357 ( .A(N2790), .B(N4745), .Y(N5425) );
  NAND2X1 gate1358 ( .A(N3813), .B(N4747), .Y(N5426) );
  NAND2X1 gate1359 ( .A(N3810), .B(N4748), .Y(N5427) );
  NAND2X1 gate1360 ( .A(N2793), .B(N4750), .Y(N5429) );
  NAND2X1 gate1361 ( .A(N3825), .B(N4752), .Y(N5430) );
  NAND2X1 gate1362 ( .A(N3822), .B(N4753), .Y(N5431) );
  NAND2X1 gate1363 ( .A(N3831), .B(N4754), .Y(N5432) );
  NAND2X1 gate1364 ( .A(N3828), .B(N4755), .Y(N5433) );
  NAND2X1 gate1365 ( .A(N2796), .B(N4775), .Y(N5451) );
  NAND2X1 gate1366 ( .A(N3864), .B(N4777), .Y(N5452) );
  NAND2X1 gate1367 ( .A(N3861), .B(N4778), .Y(N5453) );
  NAND2X1 gate1368 ( .A(N3870), .B(N4779), .Y(N5454) );
  NAND2X1 gate1369 ( .A(N3867), .B(N4780), .Y(N5455) );
  NAND2X1 gate1370 ( .A(N3888), .B(N4781), .Y(N5456) );
  NAND2X1 gate1371 ( .A(N3885), .B(N4782), .Y(N5457) );
  INVX1 gate1372 ( .A(N4303), .Y(N5469) );
  NAND2X1 gate1373 ( .A(N3589), .B(N4799), .Y(N5474) );
  NAND2X1 gate1374 ( .A(N3586), .B(N4800), .Y(N5475) );
  NAND2X1 gate1375 ( .A(N3595), .B(N4801), .Y(N5476) );
  NAND2X1 gate1376 ( .A(N3592), .B(N4802), .Y(N5477) );
  NAND2X1 gate1377 ( .A(N3798), .B(N5045), .Y(N5571) );
  NAND2X1 gate1378 ( .A(N3795), .B(N5046), .Y(N5572) );
  NAND2X1 gate1379 ( .A(N3804), .B(N5047), .Y(N5573) );
  NAND2X1 gate1380 ( .A(N3801), .B(N5048), .Y(N5574) );
  NAND2X1 gate1381 ( .A(N3837), .B(N5064), .Y(N5584) );
  NAND2X1 gate1382 ( .A(N3834), .B(N5065), .Y(N5585) );
  NAND2X1 gate1383 ( .A(N3843), .B(N5066), .Y(N5586) );
  NAND2X1 gate1384 ( .A(N3840), .B(N5067), .Y(N5587) );
  NAND2X1 gate1385 ( .A(N3876), .B(N5110), .Y(N5602) );
  NAND2X1 gate1386 ( .A(N3873), .B(N5111), .Y(N5603) );
  NAND2X1 gate1387 ( .A(N3882), .B(N5112), .Y(N5604) );
  NAND2X1 gate1388 ( .A(N3879), .B(N5113), .Y(N5605) );
  NAND2X1 gate1389 ( .A(N5324), .B(N4653), .Y(N5631) );
  NAND2X1 gate1390 ( .A(N4463), .B(N5167), .Y(N5632) );
  NAND2X1 gate1391 ( .A(N4465), .B(N5168), .Y(N5640) );
  NAND2X1 gate1392 ( .A(N4467), .B(N5169), .Y(N5654) );
  NAND2X1 gate1393 ( .A(N4469), .B(N5170), .Y(N5670) );
  NAND2X1 gate1394 ( .A(N4471), .B(N5171), .Y(N5683) );
  NAND2X1 gate1395 ( .A(N4475), .B(N5172), .Y(N5690) );
  NAND2X1 gate1396 ( .A(N4477), .B(N5173), .Y(N5697) );
  NAND2X1 gate1397 ( .A(N4479), .B(N5174), .Y(N5707) );
  NAND2X1 gate1398 ( .A(N4481), .B(N5175), .Y(N5718) );
  NAND2X1 gate1399 ( .A(N4483), .B(N5176), .Y(N5728) );
  INVX1 gate1400 ( .A(N5177), .Y(N5735) );
  NAND2X1 gate1401 ( .A(N5179), .B(N4490), .Y(N5736) );
  NAND2X1 gate1402 ( .A(N5180), .B(N5181), .Y(N5740) );
  NAND2X1 gate1403 ( .A(N5182), .B(N5183), .Y(N5744) );
  NAND2X1 gate1404 ( .A(N5184), .B(N4496), .Y(N5747) );
  NAND2X1 gate1405 ( .A(N5185), .B(N5186), .Y(N5751) );
  NAND2X1 gate1406 ( .A(N5187), .B(N5188), .Y(N5755) );
  NAND2X1 gate1407 ( .A(N5189), .B(N4502), .Y(N5758) );
  NAND2X1 gate1408 ( .A(N5190), .B(N5191), .Y(N5762) );
  NAND2X1 gate1409 ( .A(N5192), .B(N5193), .Y(N5766) );
  INVX1 gate1410 ( .A(N4803), .Y(N5769) );
  INVX1 gate1411 ( .A(N4806), .Y(N5770) );
  NAND2X1 gate1412 ( .A(N4507), .B(N5196), .Y(N5771) );
  NAND2X1 gate1413 ( .A(N4509), .B(N5197), .Y(N5778) );
  NAND2X1 gate1414 ( .A(N4511), .B(N5198), .Y(N5789) );
  NAND2X1 gate1415 ( .A(N4513), .B(N5199), .Y(N5799) );
  NAND2X1 gate1416 ( .A(N4515), .B(N5200), .Y(N5807) );
  NAND2X1 gate1417 ( .A(N4517), .B(N5201), .Y(N5821) );
  NAND2X1 gate1418 ( .A(N4519), .B(N5202), .Y(N5837) );
  NAND2X1 gate1419 ( .A(N4521), .B(N5203), .Y(N5850) );
  NAND2X1 gate1420 ( .A(N4523), .B(N5204), .Y(N5856) );
  NAND2X1 gate1421 ( .A(N4525), .B(N5205), .Y(N5863) );
  NAND2X1 gate1422 ( .A(N4527), .B(N5206), .Y(N5870) );
  NAND2X1 gate1423 ( .A(N4529), .B(N5207), .Y(N5881) );
  NAND2X1 gate1424 ( .A(N4531), .B(N5208), .Y(N5892) );
  NAND2X1 gate1425 ( .A(N4533), .B(N5209), .Y(N5898) );
  NAND2X1 gate1426 ( .A(N4535), .B(N5210), .Y(N5905) );
  NAND2X1 gate1427 ( .A(N4537), .B(N5211), .Y(N5915) );
  NAND2X1 gate1428 ( .A(N4539), .B(N5212), .Y(N5926) );
  NAND2X1 gate1429 ( .A(N4541), .B(N5213), .Y(N5936) );
  INVX1 gate1430 ( .A(N4817), .Y(N5943) );
  NAND2X1 gate1431 ( .A(N4820), .B(N1931), .Y(N5944) );
  INVX1 gate1432 ( .A(N4820), .Y(N5945) );
  NAND2X1 gate1433 ( .A(N4823), .B(N1932), .Y(N5946) );
  INVX1 gate1434 ( .A(N4823), .Y(N5947) );
  NAND2X1 gate1435 ( .A(N4826), .B(N1933), .Y(N5948) );
  INVX1 gate1436 ( .A(N4826), .Y(N5949) );
  NAND2X1 gate1437 ( .A(N4829), .B(N1934), .Y(N5950) );
  INVX1 gate1438 ( .A(N4829), .Y(N5951) );
  NAND2X1 gate1439 ( .A(N4832), .B(N1935), .Y(N5952) );
  INVX1 gate1440 ( .A(N4832), .Y(N5953) );
  NAND2X1 gate1441 ( .A(N4835), .B(N1936), .Y(N5954) );
  INVX1 gate1442 ( .A(N4835), .Y(N5955) );
  NAND2X1 gate1443 ( .A(N4838), .B(N1937), .Y(N5956) );
  INVX1 gate1444 ( .A(N4838), .Y(N5957) );
  NAND2X1 gate1445 ( .A(N4841), .B(N1938), .Y(N5958) );
  INVX1 gate1446 ( .A(N4841), .Y(N5959) );
  AND2X1 gate1447 ( .A(N2674), .B(N4769), .Y(N5960) );
  INVX1 gate1448 ( .A(N4844), .Y(N5966) );
  NAND2X1 gate1449 ( .A(N4847), .B(N1939), .Y(N5967) );
  INVX1 gate1450 ( .A(N4847), .Y(N5968) );
  NAND2X1 gate1451 ( .A(N4850), .B(N1940), .Y(N5969) );
  INVX1 gate1452 ( .A(N4850), .Y(N5970) );
  NAND2X1 gate1453 ( .A(N4853), .B(N1941), .Y(N5971) );
  INVX1 gate1454 ( .A(N4853), .Y(N5972) );
  NAND2X1 gate1455 ( .A(N4856), .B(N1942), .Y(N5973) );
  INVX1 gate1456 ( .A(N4856), .Y(N5974) );
  NAND2X1 gate1457 ( .A(N4859), .B(N1943), .Y(N5975) );
  INVX1 gate1458 ( .A(N4859), .Y(N5976) );
  NAND2X1 gate1459 ( .A(N4862), .B(N1944), .Y(N5977) );
  INVX1 gate1460 ( .A(N4862), .Y(N5978) );
  NAND2X1 gate1461 ( .A(N4865), .B(N1945), .Y(N5979) );
  INVX1 gate1462 ( .A(N4865), .Y(N5980) );
  AND2X1 gate1463 ( .A(N2674), .B(N4769), .Y(N5981) );
  NAND2X1 gate1464 ( .A(N4868), .B(N1946), .Y(N5989) );
  INVX1 gate1465 ( .A(N4868), .Y(N5990) );
  NAND2X1 gate1466 ( .A(N5283), .B(N5284), .Y(N5991) );
  NAND2X1 gate1467 ( .A(N5285), .B(N5286), .Y(N5996) );
  NAND2X1 gate1468 ( .A(N5287), .B(N5288), .Y(N6000) );
  NAND2X1 gate1469 ( .A(N5289), .B(N5290), .Y(N6003) );
  NAND2X1 gate1470 ( .A(N5291), .B(N5292), .Y(N6009) );
  NAND2X1 gate1471 ( .A(N5293), .B(N5294), .Y(N6014) );
  NAND2X1 gate1472 ( .A(N5295), .B(N5296), .Y(N6018) );
  NAND2X1 gate1473 ( .A(N5297), .B(N5298), .Y(N6021) );
  NAND2X1 gate1474 ( .A(N5299), .B(N5300), .Y(N6022) );
  INVX1 gate1475 ( .A(N4874), .Y(N6023) );
  NAND2X1 gate1476 ( .A(N4874), .B(N4629), .Y(N6024) );
  INVX1 gate1477 ( .A(N4877), .Y(N6025) );
  NAND2X1 gate1478 ( .A(N4877), .B(N4631), .Y(N6026) );
  INVX1 gate1479 ( .A(N4880), .Y(N6027) );
  NAND2X1 gate1480 ( .A(N4880), .B(N4633), .Y(N6028) );
  INVX1 gate1481 ( .A(N4883), .Y(N6029) );
  NAND2X1 gate1482 ( .A(N4883), .B(N4636), .Y(N6030) );
  INVX1 gate1483 ( .A(N4886), .Y(N6031) );
  INVX1 gate1484 ( .A(N4889), .Y(N6032) );
  INVX1 gate1485 ( .A(N4892), .Y(N6033) );
  INVX1 gate1486 ( .A(N4895), .Y(N6034) );
  INVX1 gate1487 ( .A(N4898), .Y(N6035) );
  INVX1 gate1488 ( .A(N4901), .Y(N6036) );
  INVX1 gate1489 ( .A(N4904), .Y(N6037) );
  NAND2X1 gate1490 ( .A(N4904), .B(N4642), .Y(N6038) );
  INVX1 gate1491 ( .A(N4907), .Y(N6039) );
  INVX1 gate1492 ( .A(N4910), .Y(N6040) );
  NAND2X1 gate1493 ( .A(N5314), .B(N5315), .Y(N6041) );
  NAND2X1 gate1494 ( .A(N5316), .B(N5317), .Y(N6047) );
  NAND2X1 gate1495 ( .A(N5318), .B(N5319), .Y(N6052) );
  NAND2X1 gate1496 ( .A(N5320), .B(N5321), .Y(N6056) );
  NAND2X1 gate1497 ( .A(N5322), .B(N5323), .Y(N6059) );
  NAND2X1 gate1498 ( .A(N4913), .B(N1968), .Y(N6060) );
  INVX1 gate1499 ( .A(N4913), .Y(N6061) );
  NAND2X1 gate1500 ( .A(N4916), .B(N1969), .Y(N6062) );
  INVX1 gate1501 ( .A(N4916), .Y(N6063) );
  NAND2X1 gate1502 ( .A(N4919), .B(N1970), .Y(N6064) );
  INVX1 gate1503 ( .A(N4919), .Y(N6065) );
  NAND2X1 gate1504 ( .A(N4922), .B(N1971), .Y(N6066) );
  INVX1 gate1505 ( .A(N4922), .Y(N6067) );
  NAND2X1 gate1506 ( .A(N4925), .B(N1972), .Y(N6068) );
  INVX1 gate1507 ( .A(N4925), .Y(N6069) );
  NAND2X1 gate1508 ( .A(N4928), .B(N1973), .Y(N6070) );
  INVX1 gate1509 ( .A(N4928), .Y(N6071) );
  NAND2X1 gate1510 ( .A(N4931), .B(N1974), .Y(N6072) );
  INVX1 gate1511 ( .A(N4931), .Y(N6073) );
  NAND2X1 gate1512 ( .A(N4934), .B(N1975), .Y(N6074) );
  INVX1 gate1513 ( .A(N4934), .Y(N6075) );
  NAND2X1 gate1514 ( .A(N4937), .B(N1976), .Y(N6076) );
  INVX1 gate1515 ( .A(N4937), .Y(N6077) );
  INVX1 gate1516 ( .A(N4940), .Y(N6078) );
  NAND2X1 gate1517 ( .A(N5363), .B(N4694), .Y(N6079) );
  NAND2X1 gate1518 ( .A(N5364), .B(N5365), .Y(N6083) );
  NAND2X1 gate1519 ( .A(N5366), .B(N5367), .Y(N6087) );
  INVX1 gate1520 ( .A(N4943), .Y(N6090) );
  NAND2X1 gate1521 ( .A(N4943), .B(N4699), .Y(N6091) );
  INVX1 gate1522 ( .A(N4946), .Y(N6092) );
  INVX1 gate1523 ( .A(N4949), .Y(N6093) );
  INVX1 gate1524 ( .A(N4952), .Y(N6094) );
  INVX1 gate1525 ( .A(N4955), .Y(N6095) );
  INVX1 gate1526 ( .A(N4970), .Y(N6096) );
  NAND2X1 gate1527 ( .A(N4970), .B(N4700), .Y(N6097) );
  INVX1 gate1528 ( .A(N4973), .Y(N6098) );
  INVX1 gate1529 ( .A(N4976), .Y(N6099) );
  INVX1 gate1530 ( .A(N4979), .Y(N6100) );
  INVX1 gate1531 ( .A(N4982), .Y(N6101) );
  INVX1 gate1532 ( .A(N4997), .Y(N6102) );
  NAND2X1 gate1533 ( .A(N5000), .B(N2015), .Y(N6103) );
  INVX1 gate1534 ( .A(N5000), .Y(N6104) );
  NAND2X1 gate1535 ( .A(N5003), .B(N2016), .Y(N6105) );
  INVX1 gate1536 ( .A(N5003), .Y(N6106) );
  NAND2X1 gate1537 ( .A(N5006), .B(N2017), .Y(N6107) );
  INVX1 gate1538 ( .A(N5006), .Y(N6108) );
  NAND2X1 gate1539 ( .A(N5009), .B(N2018), .Y(N6109) );
  INVX1 gate1540 ( .A(N5009), .Y(N6110) );
  NAND2X1 gate1541 ( .A(N5012), .B(N2019), .Y(N6111) );
  INVX1 gate1542 ( .A(N5012), .Y(N6112) );
  NAND2X1 gate1543 ( .A(N5015), .B(N2020), .Y(N6113) );
  INVX1 gate1544 ( .A(N5015), .Y(N6114) );
  NAND2X1 gate1545 ( .A(N5018), .B(N2021), .Y(N6115) );
  INVX1 gate1546 ( .A(N5018), .Y(N6116) );
  NAND2X1 gate1547 ( .A(N5021), .B(N2022), .Y(N6117) );
  INVX1 gate1548 ( .A(N5021), .Y(N6118) );
  NAND2X1 gate1549 ( .A(N5024), .B(N2023), .Y(N6119) );
  INVX1 gate1550 ( .A(N5024), .Y(N6120) );
  INVX1 gate1551 ( .A(N5033), .Y(N6121) );
  NAND2X1 gate1552 ( .A(N5033), .B(N4743), .Y(N6122) );
  INVX1 gate1553 ( .A(N5036), .Y(N6123) );
  INVX1 gate1554 ( .A(N5039), .Y(N6124) );
  NAND2X1 gate1555 ( .A(N5042), .B(N4744), .Y(N6125) );
  INVX1 gate1556 ( .A(N5042), .Y(N6126) );
  NAND2X1 gate1557 ( .A(N5425), .B(N4746), .Y(N6127) );
  NAND2X1 gate1558 ( .A(N5426), .B(N5427), .Y(N6131) );
  INVX1 gate1559 ( .A(N5049), .Y(N6135) );
  NAND2X1 gate1560 ( .A(N5049), .B(N4749), .Y(N6136) );
  NAND2X1 gate1561 ( .A(N5429), .B(N4751), .Y(N6137) );
  NAND2X1 gate1562 ( .A(N5430), .B(N5431), .Y(N6141) );
  NAND2X1 gate1563 ( .A(N5432), .B(N5433), .Y(N6145) );
  INVX1 gate1564 ( .A(N5068), .Y(N6148) );
  INVX1 gate1565 ( .A(N5071), .Y(N6149) );
  INVX1 gate1566 ( .A(N5074), .Y(N6150) );
  INVX1 gate1567 ( .A(N5077), .Y(N6151) );
  INVX1 gate1568 ( .A(N5080), .Y(N6152) );
  INVX1 gate1569 ( .A(N5083), .Y(N6153) );
  INVX1 gate1570 ( .A(N5086), .Y(N6154) );
  INVX1 gate1571 ( .A(N5089), .Y(N6155) );
  INVX1 gate1572 ( .A(N5092), .Y(N6156) );
  NAND2X1 gate1573 ( .A(N5092), .B(N4761), .Y(N6157) );
  INVX1 gate1574 ( .A(N5095), .Y(N6158) );
  NAND2X1 gate1575 ( .A(N5095), .B(N4763), .Y(N6159) );
  INVX1 gate1576 ( .A(N5098), .Y(N6160) );
  NAND2X1 gate1577 ( .A(N5098), .B(N4765), .Y(N6161) );
  INVX1 gate1578 ( .A(N5101), .Y(N6162) );
  INVX1 gate1579 ( .A(N5104), .Y(N6163) );
  NAND2X1 gate1580 ( .A(N5107), .B(N4768), .Y(N6164) );
  INVX1 gate1581 ( .A(N5107), .Y(N6165) );
  NAND2X1 gate1582 ( .A(N5451), .B(N4776), .Y(N6166) );
  NAND2X1 gate1583 ( .A(N5452), .B(N5453), .Y(N6170) );
  NAND2X1 gate1584 ( .A(N5454), .B(N5455), .Y(N6174) );
  NAND2X1 gate1585 ( .A(N5456), .B(N5457), .Y(N6177) );
  INVX1 gate1586 ( .A(N5114), .Y(N6181) );
  INVX1 gate1587 ( .A(N5117), .Y(N6182) );
  INVX1 gate1588 ( .A(N5120), .Y(N6183) );
  INVX1 gate1589 ( .A(N5123), .Y(N6184) );
  INVX1 gate1590 ( .A(N5138), .Y(N6185) );
  NAND2X1 gate1591 ( .A(N5138), .B(N4783), .Y(N6186) );
  INVX1 gate1592 ( .A(N5141), .Y(N6187) );
  INVX1 gate1593 ( .A(N5144), .Y(N6188) );
  INVX1 gate1594 ( .A(N5147), .Y(N6189) );
  INVX1 gate1595 ( .A(N5150), .Y(N6190) );
  INVX1 gate1596 ( .A(N4784), .Y(N6191) );
  NAND2X1 gate1597 ( .A(N4784), .B(N2230), .Y(N6192) );
  INVX1 gate1598 ( .A(N4790), .Y(N6193) );
  NAND2X1 gate1599 ( .A(N4790), .B(N2765), .Y(N6194) );
  INVX1 gate1600 ( .A(N4796), .Y(N6195) );
  NAND2X1 gate1601 ( .A(N5476), .B(N5477), .Y(N6196) );
  NAND2X1 gate1602 ( .A(N5474), .B(N5475), .Y(N6199) );
  INVX1 gate1603 ( .A(N4810), .Y(N6202) );
  INVX1 gate1604 ( .A(N4814), .Y(N6203) );
  BUFX2 gate1605 ( .A(N4769), .Y(N6204) );
  BUFX2 gate1606 ( .A(N4555), .Y(N6207) );
  BUFX2 gate1607 ( .A(N4769), .Y(N6210) );
  INVX1 gate1608 ( .A(N4871), .Y(N6213) );
  BUFX2 gate1609 ( .A(N4586), .Y(N6214) );
  NOR2X1 gate1610 ( .A(N2674), .B(N4769), .Y(N6217) );
  BUFX2 gate1611 ( .A(N4667), .Y(N6220) );
  INVX1 gate1612 ( .A(N4958), .Y(N6223) );
  INVX1 gate1613 ( .A(N4961), .Y(N6224) );
  INVX1 gate1614 ( .A(N4964), .Y(N6225) );
  INVX1 gate1615 ( .A(N4967), .Y(N6226) );
  INVX1 gate1616 ( .A(N4985), .Y(N6227) );
  INVX1 gate1617 ( .A(N4988), .Y(N6228) );
  INVX1 gate1618 ( .A(N4991), .Y(N6229) );
  INVX1 gate1619 ( .A(N4994), .Y(N6230) );
  INVX1 gate1620 ( .A(N5027), .Y(N6231) );
  BUFX2 gate1621 ( .A(N4711), .Y(N6232) );
  INVX1 gate1622 ( .A(N5030), .Y(N6235) );
  BUFX2 gate1623 ( .A(N4735), .Y(N6236) );
  INVX1 gate1624 ( .A(N5052), .Y(N6239) );
  INVX1 gate1625 ( .A(N5055), .Y(N6240) );
  INVX1 gate1626 ( .A(N5058), .Y(N6241) );
  INVX1 gate1627 ( .A(N5061), .Y(N6242) );
  NAND2X1 gate1628 ( .A(N5573), .B(N5574), .Y(N6243) );
  NAND2X1 gate1629 ( .A(N5571), .B(N5572), .Y(N6246) );
  NAND2X1 gate1630 ( .A(N5586), .B(N5587), .Y(N6249) );
  NAND2X1 gate1631 ( .A(N5584), .B(N5585), .Y(N6252) );
  INVX1 gate1632 ( .A(N5126), .Y(N6255) );
  INVX1 gate1633 ( .A(N5129), .Y(N6256) );
  INVX1 gate1634 ( .A(N5132), .Y(N6257) );
  INVX1 gate1635 ( .A(N5135), .Y(N6258) );
  INVX1 gate1636 ( .A(N5153), .Y(N6259) );
  INVX1 gate1637 ( .A(N5156), .Y(N6260) );
  INVX1 gate1638 ( .A(N5159), .Y(N6261) );
  INVX1 gate1639 ( .A(N5162), .Y(N6262) );
  NAND2X1 gate1640 ( .A(N5604), .B(N5605), .Y(N6263) );
  NAND2X1 gate1641 ( .A(N5602), .B(N5603), .Y(N6266) );
  NAND2X1 gate1642 ( .A(N1380), .B(N5945), .Y(N6540) );
  NAND2X1 gate1643 ( .A(N1383), .B(N5947), .Y(N6541) );
  NAND2X1 gate1644 ( .A(N1386), .B(N5949), .Y(N6542) );
  NAND2X1 gate1645 ( .A(N1389), .B(N5951), .Y(N6543) );
  NAND2X1 gate1646 ( .A(N1392), .B(N5953), .Y(N6544) );
  NAND2X1 gate1647 ( .A(N1395), .B(N5955), .Y(N6545) );
  NAND2X1 gate1648 ( .A(N1398), .B(N5957), .Y(N6546) );
  NAND2X1 gate1649 ( .A(N1401), .B(N5959), .Y(N6547) );
  NAND2X1 gate1650 ( .A(N1404), .B(N5968), .Y(N6555) );
  NAND2X1 gate1651 ( .A(N1407), .B(N5970), .Y(N6556) );
  NAND2X1 gate1652 ( .A(N1410), .B(N5972), .Y(N6557) );
  NAND2X1 gate1653 ( .A(N1413), .B(N5974), .Y(N6558) );
  NAND2X1 gate1654 ( .A(N1416), .B(N5976), .Y(N6559) );
  NAND2X1 gate1655 ( .A(N1419), .B(N5978), .Y(N6560) );
  NAND2X1 gate1656 ( .A(N1422), .B(N5980), .Y(N6561) );
  NAND2X1 gate1657 ( .A(N1425), .B(N5990), .Y(N6569) );
  NAND2X1 gate1658 ( .A(N3721), .B(N6023), .Y(N6594) );
  NAND2X1 gate1659 ( .A(N3724), .B(N6025), .Y(N6595) );
  NAND2X1 gate1660 ( .A(N3727), .B(N6027), .Y(N6596) );
  NAND2X1 gate1661 ( .A(N3730), .B(N6029), .Y(N6597) );
  NAND2X1 gate1662 ( .A(N4889), .B(N6031), .Y(N6598) );
  NAND2X1 gate1663 ( .A(N4886), .B(N6032), .Y(N6599) );
  NAND2X1 gate1664 ( .A(N4895), .B(N6033), .Y(N6600) );
  NAND2X1 gate1665 ( .A(N4892), .B(N6034), .Y(N6601) );
  NAND2X1 gate1666 ( .A(N4901), .B(N6035), .Y(N6602) );
  NAND2X1 gate1667 ( .A(N4898), .B(N6036), .Y(N6603) );
  NAND2X1 gate1668 ( .A(N3733), .B(N6037), .Y(N6604) );
  NAND2X1 gate1669 ( .A(N4910), .B(N6039), .Y(N6605) );
  NAND2X1 gate1670 ( .A(N4907), .B(N6040), .Y(N6606) );
  NAND2X1 gate1671 ( .A(N1434), .B(N6061), .Y(N6621) );
  NAND2X1 gate1672 ( .A(N1437), .B(N6063), .Y(N6622) );
  NAND2X1 gate1673 ( .A(N1440), .B(N6065), .Y(N6623) );
  NAND2X1 gate1674 ( .A(N1443), .B(N6067), .Y(N6624) );
  NAND2X1 gate1675 ( .A(N1446), .B(N6069), .Y(N6625) );
  NAND2X1 gate1676 ( .A(N1449), .B(N6071), .Y(N6626) );
  NAND2X1 gate1677 ( .A(N1452), .B(N6073), .Y(N6627) );
  NAND2X1 gate1678 ( .A(N1455), .B(N6075), .Y(N6628) );
  NAND2X1 gate1679 ( .A(N1458), .B(N6077), .Y(N6629) );
  NAND2X1 gate1680 ( .A(N3783), .B(N6090), .Y(N6639) );
  NAND2X1 gate1681 ( .A(N4949), .B(N6092), .Y(N6640) );
  NAND2X1 gate1682 ( .A(N4946), .B(N6093), .Y(N6641) );
  NAND2X1 gate1683 ( .A(N4955), .B(N6094), .Y(N6642) );
  NAND2X1 gate1684 ( .A(N4952), .B(N6095), .Y(N6643) );
  NAND2X1 gate1685 ( .A(N3786), .B(N6096), .Y(N6644) );
  NAND2X1 gate1686 ( .A(N4976), .B(N6098), .Y(N6645) );
  NAND2X1 gate1687 ( .A(N4973), .B(N6099), .Y(N6646) );
  NAND2X1 gate1688 ( .A(N4982), .B(N6100), .Y(N6647) );
  NAND2X1 gate1689 ( .A(N4979), .B(N6101), .Y(N6648) );
  NAND2X1 gate1690 ( .A(N1461), .B(N6104), .Y(N6649) );
  NAND2X1 gate1691 ( .A(N1464), .B(N6106), .Y(N6650) );
  NAND2X1 gate1692 ( .A(N1467), .B(N6108), .Y(N6651) );
  NAND2X1 gate1693 ( .A(N1470), .B(N6110), .Y(N6652) );
  NAND2X1 gate1694 ( .A(N1473), .B(N6112), .Y(N6653) );
  NAND2X1 gate1695 ( .A(N1476), .B(N6114), .Y(N6654) );
  NAND2X1 gate1696 ( .A(N1479), .B(N6116), .Y(N6655) );
  NAND2X1 gate1697 ( .A(N1482), .B(N6118), .Y(N6656) );
  NAND2X1 gate1698 ( .A(N1485), .B(N6120), .Y(N6657) );
  NAND2X1 gate1699 ( .A(N3789), .B(N6121), .Y(N6658) );
  NAND2X1 gate1700 ( .A(N5039), .B(N6123), .Y(N6659) );
  NAND2X1 gate1701 ( .A(N5036), .B(N6124), .Y(N6660) );
  NAND2X1 gate1702 ( .A(N3792), .B(N6126), .Y(N6661) );
  NAND2X1 gate1703 ( .A(N3816), .B(N6135), .Y(N6668) );
  NAND2X1 gate1704 ( .A(N5071), .B(N6148), .Y(N6677) );
  NAND2X1 gate1705 ( .A(N5068), .B(N6149), .Y(N6678) );
  NAND2X1 gate1706 ( .A(N5077), .B(N6150), .Y(N6679) );
  NAND2X1 gate1707 ( .A(N5074), .B(N6151), .Y(N6680) );
  NAND2X1 gate1708 ( .A(N5083), .B(N6152), .Y(N6681) );
  NAND2X1 gate1709 ( .A(N5080), .B(N6153), .Y(N6682) );
  NAND2X1 gate1710 ( .A(N5089), .B(N6154), .Y(N6683) );
  NAND2X1 gate1711 ( .A(N5086), .B(N6155), .Y(N6684) );
  NAND2X1 gate1712 ( .A(N3846), .B(N6156), .Y(N6685) );
  NAND2X1 gate1713 ( .A(N3849), .B(N6158), .Y(N6686) );
  NAND2X1 gate1714 ( .A(N3852), .B(N6160), .Y(N6687) );
  NAND2X1 gate1715 ( .A(N5104), .B(N6162), .Y(N6688) );
  NAND2X1 gate1716 ( .A(N5101), .B(N6163), .Y(N6689) );
  NAND2X1 gate1717 ( .A(N3855), .B(N6165), .Y(N6690) );
  NAND2X1 gate1718 ( .A(N5117), .B(N6181), .Y(N6702) );
  NAND2X1 gate1719 ( .A(N5114), .B(N6182), .Y(N6703) );
  NAND2X1 gate1720 ( .A(N5123), .B(N6183), .Y(N6704) );
  NAND2X1 gate1721 ( .A(N5120), .B(N6184), .Y(N6705) );
  NAND2X1 gate1722 ( .A(N3891), .B(N6185), .Y(N6706) );
  NAND2X1 gate1723 ( .A(N5144), .B(N6187), .Y(N6707) );
  NAND2X1 gate1724 ( .A(N5141), .B(N6188), .Y(N6708) );
  NAND2X1 gate1725 ( .A(N5150), .B(N6189), .Y(N6709) );
  NAND2X1 gate1726 ( .A(N5147), .B(N6190), .Y(N6710) );
  NAND2X1 gate1727 ( .A(N1708), .B(N6191), .Y(N6711) );
  NAND2X1 gate1728 ( .A(N2231), .B(N6193), .Y(N6712) );
  NAND2X1 gate1729 ( .A(N4961), .B(N6223), .Y(N6729) );
  NAND2X1 gate1730 ( .A(N4958), .B(N6224), .Y(N6730) );
  NAND2X1 gate1731 ( .A(N4967), .B(N6225), .Y(N6731) );
  NAND2X1 gate1732 ( .A(N4964), .B(N6226), .Y(N6732) );
  NAND2X1 gate1733 ( .A(N4988), .B(N6227), .Y(N6733) );
  NAND2X1 gate1734 ( .A(N4985), .B(N6228), .Y(N6734) );
  NAND2X1 gate1735 ( .A(N4994), .B(N6229), .Y(N6735) );
  NAND2X1 gate1736 ( .A(N4991), .B(N6230), .Y(N6736) );
  NAND2X1 gate1737 ( .A(N5055), .B(N6239), .Y(N6741) );
  NAND2X1 gate1738 ( .A(N5052), .B(N6240), .Y(N6742) );
  NAND2X1 gate1739 ( .A(N5061), .B(N6241), .Y(N6743) );
  NAND2X1 gate1740 ( .A(N5058), .B(N6242), .Y(N6744) );
  NAND2X1 gate1741 ( .A(N5129), .B(N6255), .Y(N6751) );
  NAND2X1 gate1742 ( .A(N5126), .B(N6256), .Y(N6752) );
  NAND2X1 gate1743 ( .A(N5135), .B(N6257), .Y(N6753) );
  NAND2X1 gate1744 ( .A(N5132), .B(N6258), .Y(N6754) );
  NAND2X1 gate1745 ( .A(N5156), .B(N6259), .Y(N6755) );
  NAND2X1 gate1746 ( .A(N5153), .B(N6260), .Y(N6756) );
  NAND2X1 gate1747 ( .A(N5162), .B(N6261), .Y(N6757) );
  NAND2X1 gate1748 ( .A(N5159), .B(N6262), .Y(N6758) );
  INVX1 gate1749 ( .A(N5892), .Y(N6761) );
  AND2X1 gate1750_1 ( .A(N5683), .B(N5670), .Y(N6762_1) );
  AND2X1 gate1750_2 ( .A(N5654), .B(N5640), .Y(N6762_2) );
  AND2X1 gate1750_3 ( .A(N5632), .B(N6762_1), .Y(N6762_3) );
  AND2X1 gate1750 ( .A(N6762_2), .B(N6762_3), .Y(N6762) );
  AND2X1 gate1751 ( .A(N5632), .B(N3097), .Y(N6766) );
  AND2X1 gate1752_1 ( .A(N5640), .B(N5632), .Y(N6767_1) );
  AND2X1 gate1752 ( .A(N3101), .B(N6767_1), .Y(N6767) );
  AND2X1 gate1753_1 ( .A(N5654), .B(N5632), .Y(N6768_1) );
  AND2X1 gate1753_2 ( .A(N3107), .B(N5640), .Y(N6768_2) );
  AND2X1 gate1753 ( .A(N6768_1), .B(N6768_2), .Y(N6768) );
  AND2X1 gate1754_1 ( .A(N5670), .B(N5654), .Y(N6769_1) );
  AND2X1 gate1754_2 ( .A(N5632), .B(N3114), .Y(N6769_2) );
  AND2X1 gate1754_3 ( .A(N5640), .B(N6769_1), .Y(N6769_3) );
  AND2X1 gate1754 ( .A(N6769_2), .B(N6769_3), .Y(N6769) );
  AND2X1 gate1755 ( .A(N5640), .B(N3101), .Y(N6770) );
  AND2X1 gate1756_1 ( .A(N5654), .B(N3107), .Y(N6771_1) );
  AND2X1 gate1756 ( .A(N5640), .B(N6771_1), .Y(N6771) );
  AND2X1 gate1757_1 ( .A(N5670), .B(N5654), .Y(N6772_1) );
  AND2X1 gate1757_2 ( .A(N3114), .B(N5640), .Y(N6772_2) );
  AND2X1 gate1757 ( .A(N6772_1), .B(N6772_2), .Y(N6772) );
  AND2X1 gate1758_1 ( .A(N5683), .B(N5654), .Y(N6773_1) );
  AND2X1 gate1758_2 ( .A(N5640), .B(N5670), .Y(N6773_2) );
  AND2X1 gate1758 ( .A(N6773_1), .B(N6773_2), .Y(N6773) );
  AND2X1 gate1759 ( .A(N5640), .B(N3101), .Y(N6774) );
  AND2X1 gate1760_1 ( .A(N5654), .B(N3107), .Y(N6775_1) );
  AND2X1 gate1760 ( .A(N5640), .B(N6775_1), .Y(N6775) );
  AND2X1 gate1761_1 ( .A(N5670), .B(N5654), .Y(N6776_1) );
  AND2X1 gate1761_2 ( .A(N3114), .B(N5640), .Y(N6776_2) );
  AND2X1 gate1761 ( .A(N6776_1), .B(N6776_2), .Y(N6776) );
  AND2X1 gate1762 ( .A(N5654), .B(N3107), .Y(N6777) );
  AND2X1 gate1763_1 ( .A(N5670), .B(N5654), .Y(N6778_1) );
  AND2X1 gate1763 ( .A(N3114), .B(N6778_1), .Y(N6778) );
  AND2X1 gate1764_1 ( .A(N5683), .B(N5654), .Y(N6779_1) );
  AND2X1 gate1764 ( .A(N5670), .B(N6779_1), .Y(N6779) );
  AND2X1 gate1765 ( .A(N5654), .B(N3107), .Y(N6780) );
  AND2X1 gate1766_1 ( .A(N5670), .B(N5654), .Y(N6781_1) );
  AND2X1 gate1766 ( .A(N3114), .B(N6781_1), .Y(N6781) );
  AND2X1 gate1767 ( .A(N5670), .B(N3114), .Y(N6782) );
  AND2X1 gate1768 ( .A(N5683), .B(N5670), .Y(N6783) );
  AND2X1 gate1769_1 ( .A(N5697), .B(N5728), .Y(N6784_1) );
  AND2X1 gate1769_2 ( .A(N5707), .B(N5690), .Y(N6784_2) );
  AND2X1 gate1769_3 ( .A(N5718), .B(N6784_1), .Y(N6784_3) );
  AND2X1 gate1769 ( .A(N6784_2), .B(N6784_3), .Y(N6784) );
  AND2X1 gate1770 ( .A(N5690), .B(N3137), .Y(N6787) );
  AND2X1 gate1771_1 ( .A(N5697), .B(N5690), .Y(N6788_1) );
  AND2X1 gate1771 ( .A(N3140), .B(N6788_1), .Y(N6788) );
  AND2X1 gate1772_1 ( .A(N5707), .B(N5690), .Y(N6789_1) );
  AND2X1 gate1772_2 ( .A(N3144), .B(N5697), .Y(N6789_2) );
  AND2X1 gate1772 ( .A(N6789_1), .B(N6789_2), .Y(N6789) );
  AND2X1 gate1773_1 ( .A(N5718), .B(N5707), .Y(N6790_1) );
  AND2X1 gate1773_2 ( .A(N5690), .B(N3149), .Y(N6790_2) );
  AND2X1 gate1773_3 ( .A(N5697), .B(N6790_1), .Y(N6790_3) );
  AND2X1 gate1773 ( .A(N6790_2), .B(N6790_3), .Y(N6790) );
  AND2X1 gate1774 ( .A(N5697), .B(N3140), .Y(N6791) );
  AND2X1 gate1775_1 ( .A(N5707), .B(N3144), .Y(N6792_1) );
  AND2X1 gate1775 ( .A(N5697), .B(N6792_1), .Y(N6792) );
  AND2X1 gate1776_1 ( .A(N5718), .B(N5707), .Y(N6793_1) );
  AND2X1 gate1776_2 ( .A(N3149), .B(N5697), .Y(N6793_2) );
  AND2X1 gate1776 ( .A(N6793_1), .B(N6793_2), .Y(N6793) );
  AND2X1 gate1777 ( .A(N3144), .B(N5707), .Y(N6794) );
  AND2X1 gate1778_1 ( .A(N5718), .B(N5707), .Y(N6795_1) );
  AND2X1 gate1778 ( .A(N3149), .B(N6795_1), .Y(N6795) );
  AND2X1 gate1779 ( .A(N5718), .B(N3149), .Y(N6796) );
  INVX1 gate1780 ( .A(N5736), .Y(N6797) );
  INVX1 gate1781 ( .A(N5740), .Y(N6800) );
  INVX1 gate1782 ( .A(N5747), .Y(N6803) );
  INVX1 gate1783 ( .A(N5751), .Y(N6806) );
  INVX1 gate1784 ( .A(N5758), .Y(N6809) );
  INVX1 gate1785 ( .A(N5762), .Y(N6812) );
  BUFX2 gate1786 ( .A(N5744), .Y(N6815) );
  BUFX2 gate1787 ( .A(N5744), .Y(N6818) );
  BUFX2 gate1788 ( .A(N5755), .Y(N6821) );
  BUFX2 gate1789 ( .A(N5755), .Y(N6824) );
  BUFX2 gate1790 ( .A(N5766), .Y(N6827) );
  BUFX2 gate1791 ( .A(N5766), .Y(N6830) );
  AND2X1 gate1792_1 ( .A(N5850), .B(N5789), .Y(N6833_1) );
  AND2X1 gate1792_2 ( .A(N5778), .B(N5771), .Y(N6833_2) );
  AND2X1 gate1792 ( .A(N6833_1), .B(N6833_2), .Y(N6833) );
  AND2X1 gate1793 ( .A(N5771), .B(N3169), .Y(N6836) );
  AND2X1 gate1794_1 ( .A(N5778), .B(N5771), .Y(N6837_1) );
  AND2X1 gate1794 ( .A(N3173), .B(N6837_1), .Y(N6837) );
  AND2X1 gate1795_1 ( .A(N5789), .B(N5771), .Y(N6838_1) );
  AND2X1 gate1795_2 ( .A(N3178), .B(N5778), .Y(N6838_2) );
  AND2X1 gate1795 ( .A(N6838_1), .B(N6838_2), .Y(N6838) );
  AND2X1 gate1796 ( .A(N5778), .B(N3173), .Y(N6839) );
  AND2X1 gate1797_1 ( .A(N5789), .B(N3178), .Y(N6840_1) );
  AND2X1 gate1797 ( .A(N5778), .B(N6840_1), .Y(N6840) );
  AND2X1 gate1798_1 ( .A(N5850), .B(N5789), .Y(N6841_1) );
  AND2X1 gate1798 ( .A(N5778), .B(N6841_1), .Y(N6841) );
  AND2X1 gate1799 ( .A(N5778), .B(N3173), .Y(N6842) );
  AND2X1 gate1800_1 ( .A(N5789), .B(N3178), .Y(N6843_1) );
  AND2X1 gate1800 ( .A(N5778), .B(N6843_1), .Y(N6843) );
  AND2X1 gate1801 ( .A(N5789), .B(N3178), .Y(N6844) );
  AND2X1 gate1802_1 ( .A(N5856), .B(N5837), .Y(N6845_1) );
  AND2X1 gate1802_2 ( .A(N5821), .B(N5807), .Y(N6845_2) );
  AND2X1 gate1802_3 ( .A(N5799), .B(N6845_1), .Y(N6845_3) );
  AND2X1 gate1802 ( .A(N6845_2), .B(N6845_3), .Y(N6845) );
  AND2X1 gate1803 ( .A(N5799), .B(N3185), .Y(N6848) );
  AND2X1 gate1804_1 ( .A(N5807), .B(N5799), .Y(N6849_1) );
  AND2X1 gate1804 ( .A(N3189), .B(N6849_1), .Y(N6849) );
  AND2X1 gate1805_1 ( .A(N5821), .B(N5799), .Y(N6850_1) );
  AND2X1 gate1805_2 ( .A(N3195), .B(N5807), .Y(N6850_2) );
  AND2X1 gate1805 ( .A(N6850_1), .B(N6850_2), .Y(N6850) );
  AND2X1 gate1806_1 ( .A(N5837), .B(N5821), .Y(N6851_1) );
  AND2X1 gate1806_2 ( .A(N5799), .B(N3202), .Y(N6851_2) );
  AND2X1 gate1806_3 ( .A(N5807), .B(N6851_1), .Y(N6851_3) );
  AND2X1 gate1806 ( .A(N6851_2), .B(N6851_3), .Y(N6851) );
  AND2X1 gate1807 ( .A(N5807), .B(N3189), .Y(N6852) );
  AND2X1 gate1808_1 ( .A(N5821), .B(N3195), .Y(N6853_1) );
  AND2X1 gate1808 ( .A(N5807), .B(N6853_1), .Y(N6853) );
  AND2X1 gate1809_1 ( .A(N5837), .B(N5821), .Y(N6854_1) );
  AND2X1 gate1809_2 ( .A(N3202), .B(N5807), .Y(N6854_2) );
  AND2X1 gate1809 ( .A(N6854_1), .B(N6854_2), .Y(N6854) );
  AND2X1 gate1810_1 ( .A(N5856), .B(N5821), .Y(N6855_1) );
  AND2X1 gate1810_2 ( .A(N5807), .B(N5837), .Y(N6855_2) );
  AND2X1 gate1810 ( .A(N6855_1), .B(N6855_2), .Y(N6855) );
  AND2X1 gate1811 ( .A(N5807), .B(N3189), .Y(N6856) );
  AND2X1 gate1812_1 ( .A(N5821), .B(N3195), .Y(N6857_1) );
  AND2X1 gate1812 ( .A(N5807), .B(N6857_1), .Y(N6857) );
  AND2X1 gate1813_1 ( .A(N5837), .B(N5821), .Y(N6858_1) );
  AND2X1 gate1813_2 ( .A(N3202), .B(N5807), .Y(N6858_2) );
  AND2X1 gate1813 ( .A(N6858_1), .B(N6858_2), .Y(N6858) );
  AND2X1 gate1814 ( .A(N5821), .B(N3195), .Y(N6859) );
  AND2X1 gate1815_1 ( .A(N5837), .B(N5821), .Y(N6860_1) );
  AND2X1 gate1815 ( .A(N3202), .B(N6860_1), .Y(N6860) );
  AND2X1 gate1816_1 ( .A(N5856), .B(N5821), .Y(N6861_1) );
  AND2X1 gate1816 ( .A(N5837), .B(N6861_1), .Y(N6861) );
  AND2X1 gate1817 ( .A(N5821), .B(N3195), .Y(N6862) );
  AND2X1 gate1818_1 ( .A(N5837), .B(N5821), .Y(N6863_1) );
  AND2X1 gate1818 ( .A(N3202), .B(N6863_1), .Y(N6863) );
  AND2X1 gate1819 ( .A(N5837), .B(N3202), .Y(N6864) );
  AND2X1 gate1820 ( .A(N5850), .B(N5789), .Y(N6865) );
  AND2X1 gate1821 ( .A(N5856), .B(N5837), .Y(N6866) );
  AND2X1 gate1822_1 ( .A(N5870), .B(N5892), .Y(N6867_1) );
  AND2X1 gate1822_2 ( .A(N5881), .B(N5863), .Y(N6867_2) );
  AND2X1 gate1822 ( .A(N6867_1), .B(N6867_2), .Y(N6867) );
  AND2X1 gate1823 ( .A(N5863), .B(N3211), .Y(N6870) );
  AND2X1 gate1824_1 ( .A(N5870), .B(N5863), .Y(N6871_1) );
  AND2X1 gate1824 ( .A(N3215), .B(N6871_1), .Y(N6871) );
  AND2X1 gate1825_1 ( .A(N5881), .B(N5863), .Y(N6872_1) );
  AND2X1 gate1825_2 ( .A(N3221), .B(N5870), .Y(N6872_2) );
  AND2X1 gate1825 ( .A(N6872_1), .B(N6872_2), .Y(N6872) );
  AND2X1 gate1826 ( .A(N5870), .B(N3215), .Y(N6873) );
  AND2X1 gate1827_1 ( .A(N5881), .B(N3221), .Y(N6874_1) );
  AND2X1 gate1827 ( .A(N5870), .B(N6874_1), .Y(N6874) );
  AND2X1 gate1828_1 ( .A(N5892), .B(N5881), .Y(N6875_1) );
  AND2X1 gate1828 ( .A(N5870), .B(N6875_1), .Y(N6875) );
  AND2X1 gate1829 ( .A(N5870), .B(N3215), .Y(N6876) );
  AND2X1 gate1830_1 ( .A(N3221), .B(N5881), .Y(N6877_1) );
  AND2X1 gate1830 ( .A(N5870), .B(N6877_1), .Y(N6877) );
  AND2X1 gate1831 ( .A(N5881), .B(N3221), .Y(N6878) );
  AND2X1 gate1832 ( .A(N5892), .B(N5881), .Y(N6879) );
  AND2X1 gate1833 ( .A(N5881), .B(N3221), .Y(N6880) );
  AND2X1 gate1834_1 ( .A(N5905), .B(N5936), .Y(N6881_1) );
  AND2X1 gate1834_2 ( .A(N5915), .B(N5898), .Y(N6881_2) );
  AND2X1 gate1834_3 ( .A(N5926), .B(N6881_1), .Y(N6881_3) );
  AND2X1 gate1834 ( .A(N6881_2), .B(N6881_3), .Y(N6881) );
  AND2X1 gate1835 ( .A(N5898), .B(N3229), .Y(N6884) );
  AND2X1 gate1836_1 ( .A(N5905), .B(N5898), .Y(N6885_1) );
  AND2X1 gate1836 ( .A(N3232), .B(N6885_1), .Y(N6885) );
  AND2X1 gate1837_1 ( .A(N5915), .B(N5898), .Y(N6886_1) );
  AND2X1 gate1837_2 ( .A(N3236), .B(N5905), .Y(N6886_2) );
  AND2X1 gate1837 ( .A(N6886_1), .B(N6886_2), .Y(N6886) );
  AND2X1 gate1838_1 ( .A(N5926), .B(N5915), .Y(N6887_1) );
  AND2X1 gate1838_2 ( .A(N5898), .B(N3241), .Y(N6887_2) );
  AND2X1 gate1838_3 ( .A(N5905), .B(N6887_1), .Y(N6887_3) );
  AND2X1 gate1838 ( .A(N6887_2), .B(N6887_3), .Y(N6887) );
  AND2X1 gate1839 ( .A(N5905), .B(N3232), .Y(N6888) );
  AND2X1 gate1840_1 ( .A(N5915), .B(N3236), .Y(N6889_1) );
  AND2X1 gate1840 ( .A(N5905), .B(N6889_1), .Y(N6889) );
  AND2X1 gate1841_1 ( .A(N5926), .B(N5915), .Y(N6890_1) );
  AND2X1 gate1841_2 ( .A(N3241), .B(N5905), .Y(N6890_2) );
  AND2X1 gate1841 ( .A(N6890_1), .B(N6890_2), .Y(N6890) );
  AND2X1 gate1842 ( .A(N3236), .B(N5915), .Y(N6891) );
  AND2X1 gate1843_1 ( .A(N5926), .B(N5915), .Y(N6892_1) );
  AND2X1 gate1843 ( .A(N3241), .B(N6892_1), .Y(N6892) );
  AND2X1 gate1844 ( .A(N5926), .B(N3241), .Y(N6893) );
  NAND2X1 gate1845 ( .A(N5944), .B(N6540), .Y(N6894) );
  NAND2X1 gate1846 ( .A(N5946), .B(N6541), .Y(N6901) );
  NAND2X1 gate1847 ( .A(N5948), .B(N6542), .Y(N6912) );
  NAND2X1 gate1848 ( .A(N5950), .B(N6543), .Y(N6923) );
  NAND2X1 gate1849 ( .A(N5952), .B(N6544), .Y(N6929) );
  NAND2X1 gate1850 ( .A(N5954), .B(N6545), .Y(N6936) );
  NAND2X1 gate1851 ( .A(N5956), .B(N6546), .Y(N6946) );
  NAND2X1 gate1852 ( .A(N5958), .B(N6547), .Y(N6957) );
  NAND2X1 gate1853 ( .A(N6204), .B(N4575), .Y(N6967) );
  INVX1 gate1854 ( .A(N6204), .Y(N6968) );
  INVX1 gate1855 ( .A(N6207), .Y(N6969) );
  NAND2X1 gate1856 ( .A(N5967), .B(N6555), .Y(N6970) );
  NAND2X1 gate1857 ( .A(N5969), .B(N6556), .Y(N6977) );
  NAND2X1 gate1858 ( .A(N5971), .B(N6557), .Y(N6988) );
  NAND2X1 gate1859 ( .A(N5973), .B(N6558), .Y(N6998) );
  NAND2X1 gate1860 ( .A(N5975), .B(N6559), .Y(N7006) );
  NAND2X1 gate1861 ( .A(N5977), .B(N6560), .Y(N7020) );
  NAND2X1 gate1862 ( .A(N5979), .B(N6561), .Y(N7036) );
  NAND2X1 gate1863 ( .A(N5989), .B(N6569), .Y(N7049) );
  NAND2X1 gate1864 ( .A(N6210), .B(N4610), .Y(N7055) );
  INVX1 gate1865 ( .A(N6210), .Y(N7056) );
  AND2X1 gate1866_1 ( .A(N6021), .B(N6000), .Y(N7057_1) );
  AND2X1 gate1866_2 ( .A(N5996), .B(N5991), .Y(N7057_2) );
  AND2X1 gate1866 ( .A(N7057_1), .B(N7057_2), .Y(N7057) );
  AND2X1 gate1867 ( .A(N5991), .B(N3362), .Y(N7060) );
  AND2X1 gate1868_1 ( .A(N5996), .B(N5991), .Y(N7061_1) );
  AND2X1 gate1868 ( .A(N3363), .B(N7061_1), .Y(N7061) );
  AND2X1 gate1869_1 ( .A(N6000), .B(N5991), .Y(N7062_1) );
  AND2X1 gate1869_2 ( .A(N3364), .B(N5996), .Y(N7062_2) );
  AND2X1 gate1869 ( .A(N7062_1), .B(N7062_2), .Y(N7062) );
  AND2X1 gate1870_1 ( .A(N6022), .B(N6018), .Y(N7063_1) );
  AND2X1 gate1870_2 ( .A(N6014), .B(N6009), .Y(N7063_2) );
  AND2X1 gate1870_3 ( .A(N6003), .B(N7063_1), .Y(N7063_3) );
  AND2X1 gate1870 ( .A(N7063_2), .B(N7063_3), .Y(N7063) );
  AND2X1 gate1871 ( .A(N6003), .B(N3366), .Y(N7064) );
  AND2X1 gate1872_1 ( .A(N6009), .B(N6003), .Y(N7065_1) );
  AND2X1 gate1872 ( .A(N3367), .B(N7065_1), .Y(N7065) );
  AND2X1 gate1873_1 ( .A(N6014), .B(N6003), .Y(N7066_1) );
  AND2X1 gate1873_2 ( .A(N3368), .B(N6009), .Y(N7066_2) );
  AND2X1 gate1873 ( .A(N7066_1), .B(N7066_2), .Y(N7066) );
  AND2X1 gate1874_1 ( .A(N6018), .B(N6014), .Y(N7067_1) );
  AND2X1 gate1874_2 ( .A(N6003), .B(N3369), .Y(N7067_2) );
  AND2X1 gate1874_3 ( .A(N6009), .B(N7067_1), .Y(N7067_3) );
  AND2X1 gate1874 ( .A(N7067_2), .B(N7067_3), .Y(N7067) );
  NAND2X1 gate1875 ( .A(N6594), .B(N6024), .Y(N7068) );
  NAND2X1 gate1876 ( .A(N6595), .B(N6026), .Y(N7073) );
  NAND2X1 gate1877 ( .A(N6596), .B(N6028), .Y(N7077) );
  NAND2X1 gate1878 ( .A(N6597), .B(N6030), .Y(N7080) );
  NAND2X1 gate1879 ( .A(N6598), .B(N6599), .Y(N7086) );
  NAND2X1 gate1880 ( .A(N6600), .B(N6601), .Y(N7091) );
  NAND2X1 gate1881 ( .A(N6602), .B(N6603), .Y(N7095) );
  NAND2X1 gate1882 ( .A(N6604), .B(N6038), .Y(N7098) );
  NAND2X1 gate1883 ( .A(N6605), .B(N6606), .Y(N7099) );
  AND2X1 gate1884_1 ( .A(N6059), .B(N6056), .Y(N7100_1) );
  AND2X1 gate1884_2 ( .A(N6052), .B(N6047), .Y(N7100_2) );
  AND2X1 gate1884_3 ( .A(N6041), .B(N7100_1), .Y(N7100_3) );
  AND2X1 gate1884 ( .A(N7100_2), .B(N7100_3), .Y(N7100) );
  AND2X1 gate1885 ( .A(N6041), .B(N3371), .Y(N7103) );
  AND2X1 gate1886_1 ( .A(N6047), .B(N6041), .Y(N7104_1) );
  AND2X1 gate1886 ( .A(N3372), .B(N7104_1), .Y(N7104) );
  AND2X1 gate1887_1 ( .A(N6052), .B(N6041), .Y(N7105_1) );
  AND2X1 gate1887_2 ( .A(N3373), .B(N6047), .Y(N7105_2) );
  AND2X1 gate1887 ( .A(N7105_1), .B(N7105_2), .Y(N7105) );
  AND2X1 gate1888_1 ( .A(N6056), .B(N6052), .Y(N7106_1) );
  AND2X1 gate1888_2 ( .A(N6041), .B(N3374), .Y(N7106_2) );
  AND2X1 gate1888_3 ( .A(N6047), .B(N7106_1), .Y(N7106_3) );
  AND2X1 gate1888 ( .A(N7106_2), .B(N7106_3), .Y(N7106) );
  NAND2X1 gate1889 ( .A(N6060), .B(N6621), .Y(N7107) );
  NAND2X1 gate1890 ( .A(N6062), .B(N6622), .Y(N7114) );
  NAND2X1 gate1891 ( .A(N6064), .B(N6623), .Y(N7125) );
  NAND2X1 gate1892 ( .A(N6066), .B(N6624), .Y(N7136) );
  NAND2X1 gate1893 ( .A(N6068), .B(N6625), .Y(N7142) );
  NAND2X1 gate1894 ( .A(N6070), .B(N6626), .Y(N7149) );
  NAND2X1 gate1895 ( .A(N6072), .B(N6627), .Y(N7159) );
  NAND2X1 gate1896 ( .A(N6074), .B(N6628), .Y(N7170) );
  NAND2X1 gate1897 ( .A(N6076), .B(N6629), .Y(N7180) );
  INVX1 gate1898 ( .A(N6220), .Y(N7187) );
  INVX1 gate1899 ( .A(N6079), .Y(N7188) );
  INVX1 gate1900 ( .A(N6083), .Y(N7191) );
  NAND2X1 gate1901 ( .A(N6639), .B(N6091), .Y(N7194) );
  NAND2X1 gate1902 ( .A(N6640), .B(N6641), .Y(N7198) );
  NAND2X1 gate1903 ( .A(N6642), .B(N6643), .Y(N7202) );
  NAND2X1 gate1904 ( .A(N6644), .B(N6097), .Y(N7205) );
  NAND2X1 gate1905 ( .A(N6645), .B(N6646), .Y(N7209) );
  NAND2X1 gate1906 ( .A(N6647), .B(N6648), .Y(N7213) );
  BUFX2 gate1907 ( .A(N6087), .Y(N7216) );
  BUFX2 gate1908 ( .A(N6087), .Y(N7219) );
  NAND2X1 gate1909 ( .A(N6103), .B(N6649), .Y(N7222) );
  NAND2X1 gate1910 ( .A(N6105), .B(N6650), .Y(N7229) );
  NAND2X1 gate1911 ( .A(N6107), .B(N6651), .Y(N7240) );
  NAND2X1 gate1912 ( .A(N6109), .B(N6652), .Y(N7250) );
  NAND2X1 gate1913 ( .A(N6111), .B(N6653), .Y(N7258) );
  NAND2X1 gate1914 ( .A(N6113), .B(N6654), .Y(N7272) );
  NAND2X1 gate1915 ( .A(N6115), .B(N6655), .Y(N7288) );
  NAND2X1 gate1916 ( .A(N6117), .B(N6656), .Y(N7301) );
  NAND2X1 gate1917 ( .A(N6119), .B(N6657), .Y(N7307) );
  NAND2X1 gate1918 ( .A(N6658), .B(N6122), .Y(N7314) );
  NAND2X1 gate1919 ( .A(N6659), .B(N6660), .Y(N7318) );
  NAND2X1 gate1920 ( .A(N6125), .B(N6661), .Y(N7322) );
  INVX1 gate1921 ( .A(N6127), .Y(N7325) );
  INVX1 gate1922 ( .A(N6131), .Y(N7328) );
  NAND2X1 gate1923 ( .A(N6668), .B(N6136), .Y(N7331) );
  INVX1 gate1924 ( .A(N6137), .Y(N7334) );
  INVX1 gate1925 ( .A(N6141), .Y(N7337) );
  BUFX2 gate1926 ( .A(N6145), .Y(N7340) );
  BUFX2 gate1927 ( .A(N6145), .Y(N7343) );
  NAND2X1 gate1928 ( .A(N6677), .B(N6678), .Y(N7346) );
  NAND2X1 gate1929 ( .A(N6679), .B(N6680), .Y(N7351) );
  NAND2X1 gate1930 ( .A(N6681), .B(N6682), .Y(N7355) );
  NAND2X1 gate1931 ( .A(N6683), .B(N6684), .Y(N7358) );
  NAND2X1 gate1932 ( .A(N6685), .B(N6157), .Y(N7364) );
  NAND2X1 gate1933 ( .A(N6686), .B(N6159), .Y(N7369) );
  NAND2X1 gate1934 ( .A(N6687), .B(N6161), .Y(N7373) );
  NAND2X1 gate1935 ( .A(N6688), .B(N6689), .Y(N7376) );
  NAND2X1 gate1936 ( .A(N6164), .B(N6690), .Y(N7377) );
  INVX1 gate1937 ( .A(N6166), .Y(N7378) );
  INVX1 gate1938 ( .A(N6170), .Y(N7381) );
  INVX1 gate1939 ( .A(N6177), .Y(N7384) );
  NAND2X1 gate1940 ( .A(N6702), .B(N6703), .Y(N7387) );
  NAND2X1 gate1941 ( .A(N6704), .B(N6705), .Y(N7391) );
  NAND2X1 gate1942 ( .A(N6706), .B(N6186), .Y(N7394) );
  NAND2X1 gate1943 ( .A(N6707), .B(N6708), .Y(N7398) );
  NAND2X1 gate1944 ( .A(N6709), .B(N6710), .Y(N7402) );
  BUFX2 gate1945 ( .A(N6174), .Y(N7405) );
  BUFX2 gate1946 ( .A(N6174), .Y(N7408) );
  BUFX2 gate1947 ( .A(N5936), .Y(N7411) );
  BUFX2 gate1948 ( .A(N5898), .Y(N7414) );
  BUFX2 gate1949 ( .A(N5905), .Y(N7417) );
  BUFX2 gate1950 ( .A(N5915), .Y(N7420) );
  BUFX2 gate1951 ( .A(N5926), .Y(N7423) );
  BUFX2 gate1952 ( .A(N5728), .Y(N7426) );
  BUFX2 gate1953 ( .A(N5690), .Y(N7429) );
  BUFX2 gate1954 ( .A(N5697), .Y(N7432) );
  BUFX2 gate1955 ( .A(N5707), .Y(N7435) );
  BUFX2 gate1956 ( .A(N5718), .Y(N7438) );
  NAND2X1 gate1957 ( .A(N6192), .B(N6711), .Y(N7441) );
  NAND2X1 gate1958 ( .A(N6194), .B(N6712), .Y(N7444) );
  BUFX2 gate1959 ( .A(N5683), .Y(N7447) );
  BUFX2 gate1960 ( .A(N5670), .Y(N7450) );
  BUFX2 gate1961 ( .A(N5632), .Y(N7453) );
  BUFX2 gate1962 ( .A(N5654), .Y(N7456) );
  BUFX2 gate1963 ( .A(N5640), .Y(N7459) );
  BUFX2 gate1964 ( .A(N5640), .Y(N7462) );
  BUFX2 gate1965 ( .A(N5683), .Y(N7465) );
  BUFX2 gate1966 ( .A(N5670), .Y(N7468) );
  BUFX2 gate1967 ( .A(N5632), .Y(N7471) );
  BUFX2 gate1968 ( .A(N5654), .Y(N7474) );
  INVX1 gate1969 ( .A(N6196), .Y(N7477) );
  INVX1 gate1970 ( .A(N6199), .Y(N7478) );
  BUFX2 gate1971 ( .A(N5850), .Y(N7479) );
  BUFX2 gate1972 ( .A(N5789), .Y(N7482) );
  BUFX2 gate1973 ( .A(N5771), .Y(N7485) );
  BUFX2 gate1974 ( .A(N5778), .Y(N7488) );
  BUFX2 gate1975 ( .A(N5850), .Y(N7491) );
  BUFX2 gate1976 ( .A(N5789), .Y(N7494) );
  BUFX2 gate1977 ( .A(N5771), .Y(N7497) );
  BUFX2 gate1978 ( .A(N5778), .Y(N7500) );
  BUFX2 gate1979 ( .A(N5856), .Y(N7503) );
  BUFX2 gate1980 ( .A(N5837), .Y(N7506) );
  BUFX2 gate1981 ( .A(N5799), .Y(N7509) );
  BUFX2 gate1982 ( .A(N5821), .Y(N7512) );
  BUFX2 gate1983 ( .A(N5807), .Y(N7515) );
  BUFX2 gate1984 ( .A(N5807), .Y(N7518) );
  BUFX2 gate1985 ( .A(N5856), .Y(N7521) );
  BUFX2 gate1986 ( .A(N5837), .Y(N7524) );
  BUFX2 gate1987 ( .A(N5799), .Y(N7527) );
  BUFX2 gate1988 ( .A(N5821), .Y(N7530) );
  BUFX2 gate1989 ( .A(N5863), .Y(N7533) );
  BUFX2 gate1990 ( .A(N5863), .Y(N7536) );
  BUFX2 gate1991 ( .A(N5870), .Y(N7539) );
  BUFX2 gate1992 ( .A(N5870), .Y(N7542) );
  BUFX2 gate1993 ( .A(N5881), .Y(N7545) );
  BUFX2 gate1994 ( .A(N5881), .Y(N7548) );
  INVX1 gate1995 ( .A(N6214), .Y(N7551) );
  INVX1 gate1996 ( .A(N6217), .Y(N7552) );
  BUFX2 gate1997 ( .A(N5981), .Y(N7553) );
  INVX1 gate1998 ( .A(N6249), .Y(N7556) );
  INVX1 gate1999 ( .A(N6252), .Y(N7557) );
  INVX1 gate2000 ( .A(N6243), .Y(N7558) );
  INVX1 gate2001 ( .A(N6246), .Y(N7559) );
  NAND2X1 gate2002 ( .A(N6731), .B(N6732), .Y(N7560) );
  NAND2X1 gate2003 ( .A(N6729), .B(N6730), .Y(N7563) );
  NAND2X1 gate2004 ( .A(N6735), .B(N6736), .Y(N7566) );
  NAND2X1 gate2005 ( .A(N6733), .B(N6734), .Y(N7569) );
  INVX1 gate2006 ( .A(N6232), .Y(N7572) );
  INVX1 gate2007 ( .A(N6236), .Y(N7573) );
  NAND2X1 gate2008 ( .A(N6743), .B(N6744), .Y(N7574) );
  NAND2X1 gate2009 ( .A(N6741), .B(N6742), .Y(N7577) );
  INVX1 gate2010 ( .A(N6263), .Y(N7580) );
  INVX1 gate2011 ( .A(N6266), .Y(N7581) );
  NAND2X1 gate2012 ( .A(N6753), .B(N6754), .Y(N7582) );
  NAND2X1 gate2013 ( .A(N6751), .B(N6752), .Y(N7585) );
  NAND2X1 gate2014 ( .A(N6757), .B(N6758), .Y(N7588) );
  NAND2X1 gate2015 ( .A(N6755), .B(N6756), .Y(N7591) );
  OR2X1 gate2016_1 ( .A(N3096), .B(N6766), .Y(N7609_1) );
  OR2X1 gate2016_2 ( .A(N6767), .B(N6768), .Y(N7609_2) );
  OR2X1 gate2016_3 ( .A(N6769), .B(N7609_1), .Y(N7609_3) );
  OR2X1 gate2016 ( .A(N7609_2), .B(N7609_3), .Y(N7609) );
  OR2X1 gate2017 ( .A(N3107), .B(N6782), .Y(N7613) );
  OR2X1 gate2018_1 ( .A(N3136), .B(N6787), .Y(N7620_1) );
  OR2X1 gate2018_2 ( .A(N6788), .B(N6789), .Y(N7620_2) );
  OR2X1 gate2018_3 ( .A(N6790), .B(N7620_1), .Y(N7620_3) );
  OR2X1 gate2018 ( .A(N7620_2), .B(N7620_3), .Y(N7620) );
  OR2X1 gate2019_1 ( .A(N3168), .B(N6836), .Y(N7649_1) );
  OR2X1 gate2019_2 ( .A(N6837), .B(N6838), .Y(N7649_2) );
  OR2X1 gate2019 ( .A(N7649_1), .B(N7649_2), .Y(N7649) );
  OR2X1 gate2020 ( .A(N3173), .B(N6844), .Y(N7650) );
  OR2X1 gate2021_1 ( .A(N3184), .B(N6848), .Y(N7655_1) );
  OR2X1 gate2021_2 ( .A(N6849), .B(N6850), .Y(N7655_2) );
  OR2X1 gate2021_3 ( .A(N6851), .B(N7655_1), .Y(N7655_3) );
  OR2X1 gate2021 ( .A(N7655_2), .B(N7655_3), .Y(N7655) );
  OR2X1 gate2022 ( .A(N3195), .B(N6864), .Y(N7659) );
  OR2X1 gate2023_1 ( .A(N3210), .B(N6870), .Y(N7668_1) );
  OR2X1 gate2023_2 ( .A(N6871), .B(N6872), .Y(N7668_2) );
  OR2X1 gate2023 ( .A(N7668_1), .B(N7668_2), .Y(N7668) );
  OR2X1 gate2024_1 ( .A(N3228), .B(N6884), .Y(N7671_1) );
  OR2X1 gate2024_2 ( .A(N6885), .B(N6886), .Y(N7671_2) );
  OR2X1 gate2024_3 ( .A(N6887), .B(N7671_1), .Y(N7671_3) );
  OR2X1 gate2024 ( .A(N7671_2), .B(N7671_3), .Y(N7671) );
  NAND2X1 gate2025 ( .A(N3661), .B(N6968), .Y(N7744) );
  NAND2X1 gate2026 ( .A(N3664), .B(N7056), .Y(N7822) );
  OR2X1 gate2027_1 ( .A(N3361), .B(N7060), .Y(N7825_1) );
  OR2X1 gate2027_2 ( .A(N7061), .B(N7062), .Y(N7825_2) );
  OR2X1 gate2027 ( .A(N7825_1), .B(N7825_2), .Y(N7825) );
  OR2X1 gate2028_1 ( .A(N3365), .B(N7064), .Y(N7826_1) );
  OR2X1 gate2028_2 ( .A(N7065), .B(N7066), .Y(N7826_2) );
  OR2X1 gate2028_3 ( .A(N7067), .B(N7826_1), .Y(N7826_3) );
  OR2X1 gate2028 ( .A(N7826_2), .B(N7826_3), .Y(N7826) );
  OR2X1 gate2029_1 ( .A(N3370), .B(N7103), .Y(N7852_1) );
  OR2X1 gate2029_2 ( .A(N7104), .B(N7105), .Y(N7852_2) );
  OR2X1 gate2029_3 ( .A(N7106), .B(N7852_1), .Y(N7852_3) );
  OR2X1 gate2029 ( .A(N7852_2), .B(N7852_3), .Y(N7852) );
  OR2X1 gate2030_1 ( .A(N3101), .B(N6777), .Y(N8114_1) );
  OR2X1 gate2030_2 ( .A(N6778), .B(N6779), .Y(N8114_2) );
  OR2X1 gate2030 ( .A(N8114_1), .B(N8114_2), .Y(N8114) );
  OR2X1 gate2031_1 ( .A(N3097), .B(N6770), .Y(N8117_1) );
  OR2X1 gate2031_2 ( .A(N6771), .B(N6772), .Y(N8117_2) );
  OR2X1 gate2031_3 ( .A(N6773), .B(N8117_1), .Y(N8117_3) );
  OR2X1 gate2031 ( .A(N8117_2), .B(N8117_3), .Y(N8117) );
  NOR3X1 gate2032 ( .A(N3101), .B(N6780), .C(N6781), .Y(N8131) );
  NOR2X1 gate2033_1 ( .A(N3097), .B(N6774), .Y(N8134_1) );
  NOR2X1 gate2033_2 ( .A(N6775), .B(N6776), .Y(N8134_2) );
  NOR2X1 gate2033 ( .A(N8134_1), .B(N8134_2), .Y(N8134) );
  NAND2X1 gate2034 ( .A(N6199), .B(N7477), .Y(N8144) );
  NAND2X1 gate2035 ( .A(N6196), .B(N7478), .Y(N8145) );
  OR2X1 gate2036_1 ( .A(N3169), .B(N6839), .Y(N8146_1) );
  OR2X1 gate2036_2 ( .A(N6840), .B(N6841), .Y(N8146_2) );
  OR2X1 gate2036 ( .A(N8146_1), .B(N8146_2), .Y(N8146) );
  NOR3X1 gate2037 ( .A(N3169), .B(N6842), .C(N6843), .Y(N8156) );
  OR2X1 gate2038_1 ( .A(N3189), .B(N6859), .Y(N8166_1) );
  OR2X1 gate2038_2 ( .A(N6860), .B(N6861), .Y(N8166_2) );
  OR2X1 gate2038 ( .A(N8166_1), .B(N8166_2), .Y(N8166) );
  OR2X1 gate2039_1 ( .A(N3185), .B(N6852), .Y(N8169_1) );
  OR2X1 gate2039_2 ( .A(N6853), .B(N6854), .Y(N8169_2) );
  OR2X1 gate2039_3 ( .A(N6855), .B(N8169_1), .Y(N8169_3) );
  OR2X1 gate2039 ( .A(N8169_2), .B(N8169_3), .Y(N8169) );
  NOR3X1 gate2040 ( .A(N3189), .B(N6862), .C(N6863), .Y(N8183) );
  NOR2X1 gate2041_1 ( .A(N3185), .B(N6856), .Y(N8186_1) );
  NOR2X1 gate2041_2 ( .A(N6857), .B(N6858), .Y(N8186_2) );
  NOR2X1 gate2041 ( .A(N8186_1), .B(N8186_2), .Y(N8186) );
  OR2X1 gate2042_1 ( .A(N3211), .B(N6873), .Y(N8196_1) );
  OR2X1 gate2042_2 ( .A(N6874), .B(N6875), .Y(N8196_2) );
  OR2X1 gate2042 ( .A(N8196_1), .B(N8196_2), .Y(N8196) );
  NOR3X1 gate2043 ( .A(N3211), .B(N6876), .C(N6877), .Y(N8200) );
  OR2X1 gate2044_1 ( .A(N3215), .B(N6878), .Y(N8204_1) );
  OR2X1 gate2044 ( .A(N6879), .B(N8204_1), .Y(N8204) );
  NOR2X1 gate2045 ( .A(N3215), .B(N6880), .Y(N8208) );
  NAND2X1 gate2046 ( .A(N6252), .B(N7556), .Y(N8216) );
  NAND2X1 gate2047 ( .A(N6249), .B(N7557), .Y(N8217) );
  NAND2X1 gate2048 ( .A(N6246), .B(N7558), .Y(N8218) );
  NAND2X1 gate2049 ( .A(N6243), .B(N7559), .Y(N8219) );
  NAND2X1 gate2050 ( .A(N6266), .B(N7580), .Y(N8232) );
  NAND2X1 gate2051 ( .A(N6263), .B(N7581), .Y(N8233) );
  INVX1 gate2052 ( .A(N7411), .Y(N8242) );
  INVX1 gate2053 ( .A(N7414), .Y(N8243) );
  INVX1 gate2054 ( .A(N7417), .Y(N8244) );
  INVX1 gate2055 ( .A(N7420), .Y(N8245) );
  INVX1 gate2056 ( .A(N7423), .Y(N8246) );
  INVX1 gate2057 ( .A(N7426), .Y(N8247) );
  INVX1 gate2058 ( .A(N7429), .Y(N8248) );
  INVX1 gate2059 ( .A(N7432), .Y(N8249) );
  INVX1 gate2060 ( .A(N7435), .Y(N8250) );
  INVX1 gate2061 ( .A(N7438), .Y(N8251) );
  INVX1 gate2062 ( .A(N7136), .Y(N8252) );
  INVX1 gate2063 ( .A(N6923), .Y(N8253) );
  INVX1 gate2064 ( .A(N6762), .Y(N8254) );
  INVX1 gate2065 ( .A(N7459), .Y(N8260) );
  INVX1 gate2066 ( .A(N7462), .Y(N8261) );
  AND2X1 gate2067 ( .A(N3122), .B(N6762), .Y(N8262) );
  AND2X1 gate2068 ( .A(N3155), .B(N6784), .Y(N8269) );
  INVX1 gate2069 ( .A(N6815), .Y(N8274) );
  INVX1 gate2070 ( .A(N6818), .Y(N8275) );
  INVX1 gate2071 ( .A(N6821), .Y(N8276) );
  INVX1 gate2072 ( .A(N6824), .Y(N8277) );
  INVX1 gate2073 ( .A(N6827), .Y(N8278) );
  INVX1 gate2074 ( .A(N6830), .Y(N8279) );
  AND2X1 gate2075_1 ( .A(N5740), .B(N5736), .Y(N8280_1) );
  AND2X1 gate2075 ( .A(N6815), .B(N8280_1), .Y(N8280) );
  AND2X1 gate2076_1 ( .A(N6800), .B(N6797), .Y(N8281_1) );
  AND2X1 gate2076 ( .A(N6818), .B(N8281_1), .Y(N8281) );
  AND2X1 gate2077_1 ( .A(N5751), .B(N5747), .Y(N8282_1) );
  AND2X1 gate2077 ( .A(N6821), .B(N8282_1), .Y(N8282) );
  AND2X1 gate2078_1 ( .A(N6806), .B(N6803), .Y(N8283_1) );
  AND2X1 gate2078 ( .A(N6824), .B(N8283_1), .Y(N8283) );
  AND2X1 gate2079_1 ( .A(N5762), .B(N5758), .Y(N8284_1) );
  AND2X1 gate2079 ( .A(N6827), .B(N8284_1), .Y(N8284) );
  AND2X1 gate2080_1 ( .A(N6812), .B(N6809), .Y(N8285_1) );
  AND2X1 gate2080 ( .A(N6830), .B(N8285_1), .Y(N8285) );
  INVX1 gate2081 ( .A(N6845), .Y(N8288) );
  INVX1 gate2082 ( .A(N7488), .Y(N8294) );
  INVX1 gate2083 ( .A(N7500), .Y(N8295) );
  INVX1 gate2084 ( .A(N7515), .Y(N8296) );
  INVX1 gate2085 ( .A(N7518), .Y(N8297) );
  AND2X1 gate2086 ( .A(N6833), .B(N6845), .Y(N8298) );
  AND2X1 gate2087 ( .A(N6867), .B(N6881), .Y(N8307) );
  INVX1 gate2088 ( .A(N7533), .Y(N8315) );
  INVX1 gate2089 ( .A(N7536), .Y(N8317) );
  INVX1 gate2090 ( .A(N7539), .Y(N8319) );
  INVX1 gate2091 ( .A(N7542), .Y(N8321) );
  NAND2X1 gate2092 ( .A(N7545), .B(N4543), .Y(N8322) );
  INVX1 gate2093 ( .A(N7545), .Y(N8323) );
  NAND2X1 gate2094 ( .A(N7548), .B(N5943), .Y(N8324) );
  INVX1 gate2095 ( .A(N7548), .Y(N8325) );
  NAND2X1 gate2096 ( .A(N6967), .B(N7744), .Y(N8326) );
  AND2X1 gate2097_1 ( .A(N6901), .B(N6923), .Y(N8333_1) );
  AND2X1 gate2097_2 ( .A(N6912), .B(N6894), .Y(N8333_2) );
  AND2X1 gate2097 ( .A(N8333_1), .B(N8333_2), .Y(N8333) );
  AND2X1 gate2098 ( .A(N6894), .B(N4545), .Y(N8337) );
  AND2X1 gate2099_1 ( .A(N6901), .B(N6894), .Y(N8338_1) );
  AND2X1 gate2099 ( .A(N4549), .B(N8338_1), .Y(N8338) );
  AND2X1 gate2100_1 ( .A(N6912), .B(N6894), .Y(N8339_1) );
  AND2X1 gate2100_2 ( .A(N4555), .B(N6901), .Y(N8339_2) );
  AND2X1 gate2100 ( .A(N8339_1), .B(N8339_2), .Y(N8339) );
  AND2X1 gate2101 ( .A(N6901), .B(N4549), .Y(N8340) );
  AND2X1 gate2102_1 ( .A(N6912), .B(N4555), .Y(N8341_1) );
  AND2X1 gate2102 ( .A(N6901), .B(N8341_1), .Y(N8341) );
  AND2X1 gate2103_1 ( .A(N6923), .B(N6912), .Y(N8342_1) );
  AND2X1 gate2103 ( .A(N6901), .B(N8342_1), .Y(N8342) );
  AND2X1 gate2104 ( .A(N6901), .B(N4549), .Y(N8343) );
  AND2X1 gate2105_1 ( .A(N4555), .B(N6912), .Y(N8344_1) );
  AND2X1 gate2105 ( .A(N6901), .B(N8344_1), .Y(N8344) );
  AND2X1 gate2106 ( .A(N6912), .B(N4555), .Y(N8345) );
  AND2X1 gate2107 ( .A(N6923), .B(N6912), .Y(N8346) );
  AND2X1 gate2108 ( .A(N6912), .B(N4555), .Y(N8347) );
  AND2X1 gate2109 ( .A(N6929), .B(N4563), .Y(N8348) );
  AND2X1 gate2110_1 ( .A(N6936), .B(N6929), .Y(N8349_1) );
  AND2X1 gate2110 ( .A(N4566), .B(N8349_1), .Y(N8349) );
  AND2X1 gate2111_1 ( .A(N6946), .B(N6929), .Y(N8350_1) );
  AND2X1 gate2111_2 ( .A(N4570), .B(N6936), .Y(N8350_2) );
  AND2X1 gate2111 ( .A(N8350_1), .B(N8350_2), .Y(N8350) );
  AND2X1 gate2112_1 ( .A(N6957), .B(N6946), .Y(N8351_1) );
  AND2X1 gate2112_2 ( .A(N6929), .B(N5960), .Y(N8351_2) );
  AND2X1 gate2112_3 ( .A(N6936), .B(N8351_1), .Y(N8351_3) );
  AND2X1 gate2112 ( .A(N8351_2), .B(N8351_3), .Y(N8351) );
  AND2X1 gate2113 ( .A(N6936), .B(N4566), .Y(N8352) );
  AND2X1 gate2114_1 ( .A(N6946), .B(N4570), .Y(N8353_1) );
  AND2X1 gate2114 ( .A(N6936), .B(N8353_1), .Y(N8353) );
  AND2X1 gate2115_1 ( .A(N6957), .B(N6946), .Y(N8354_1) );
  AND2X1 gate2115_2 ( .A(N5960), .B(N6936), .Y(N8354_2) );
  AND2X1 gate2115 ( .A(N8354_1), .B(N8354_2), .Y(N8354) );
  AND2X1 gate2116 ( .A(N4570), .B(N6946), .Y(N8355) );
  AND2X1 gate2117_1 ( .A(N6957), .B(N6946), .Y(N8356_1) );
  AND2X1 gate2117 ( .A(N5960), .B(N8356_1), .Y(N8356) );
  AND2X1 gate2118 ( .A(N6957), .B(N5960), .Y(N8357) );
  NAND2X1 gate2119 ( .A(N7055), .B(N7822), .Y(N8358) );
  AND2X1 gate2120_1 ( .A(N7049), .B(N6988), .Y(N8365_1) );
  AND2X1 gate2120_2 ( .A(N6977), .B(N6970), .Y(N8365_2) );
  AND2X1 gate2120 ( .A(N8365_1), .B(N8365_2), .Y(N8365) );
  AND2X1 gate2121 ( .A(N6970), .B(N4577), .Y(N8369) );
  AND2X1 gate2122_1 ( .A(N6977), .B(N6970), .Y(N8370_1) );
  AND2X1 gate2122 ( .A(N4581), .B(N8370_1), .Y(N8370) );
  AND2X1 gate2123_1 ( .A(N6988), .B(N6970), .Y(N8371_1) );
  AND2X1 gate2123_2 ( .A(N4586), .B(N6977), .Y(N8371_2) );
  AND2X1 gate2123 ( .A(N8371_1), .B(N8371_2), .Y(N8371) );
  AND2X1 gate2124 ( .A(N6977), .B(N4581), .Y(N8372) );
  AND2X1 gate2125_1 ( .A(N6988), .B(N4586), .Y(N8373_1) );
  AND2X1 gate2125 ( .A(N6977), .B(N8373_1), .Y(N8373) );
  AND2X1 gate2126_1 ( .A(N7049), .B(N6988), .Y(N8374_1) );
  AND2X1 gate2126 ( .A(N6977), .B(N8374_1), .Y(N8374) );
  AND2X1 gate2127 ( .A(N6977), .B(N4581), .Y(N8375) );
  AND2X1 gate2128_1 ( .A(N6988), .B(N4586), .Y(N8376_1) );
  AND2X1 gate2128 ( .A(N6977), .B(N8376_1), .Y(N8376) );
  AND2X1 gate2129 ( .A(N6988), .B(N4586), .Y(N8377) );
  AND2X1 gate2130 ( .A(N6998), .B(N4593), .Y(N8378) );
  AND2X1 gate2131_1 ( .A(N7006), .B(N6998), .Y(N8379_1) );
  AND2X1 gate2131 ( .A(N4597), .B(N8379_1), .Y(N8379) );
  AND2X1 gate2132_1 ( .A(N7020), .B(N6998), .Y(N8380_1) );
  AND2X1 gate2132_2 ( .A(N4603), .B(N7006), .Y(N8380_2) );
  AND2X1 gate2132 ( .A(N8380_1), .B(N8380_2), .Y(N8380) );
  AND2X1 gate2133_1 ( .A(N7036), .B(N7020), .Y(N8381_1) );
  AND2X1 gate2133_2 ( .A(N6998), .B(N5981), .Y(N8381_2) );
  AND2X1 gate2133_3 ( .A(N7006), .B(N8381_1), .Y(N8381_3) );
  AND2X1 gate2133 ( .A(N8381_2), .B(N8381_3), .Y(N8381) );
  AND2X1 gate2134 ( .A(N7006), .B(N4597), .Y(N8382) );
  AND2X1 gate2135_1 ( .A(N7020), .B(N4603), .Y(N8383_1) );
  AND2X1 gate2135 ( .A(N7006), .B(N8383_1), .Y(N8383) );
  AND2X1 gate2136_1 ( .A(N7036), .B(N7020), .Y(N8384_1) );
  AND2X1 gate2136_2 ( .A(N5981), .B(N7006), .Y(N8384_2) );
  AND2X1 gate2136 ( .A(N8384_1), .B(N8384_2), .Y(N8384) );
  AND2X1 gate2137 ( .A(N7006), .B(N4597), .Y(N8385) );
  AND2X1 gate2138_1 ( .A(N7020), .B(N4603), .Y(N8386_1) );
  AND2X1 gate2138 ( .A(N7006), .B(N8386_1), .Y(N8386) );
  AND2X1 gate2139_1 ( .A(N7036), .B(N7020), .Y(N8387_1) );
  AND2X1 gate2139_2 ( .A(N5981), .B(N7006), .Y(N8387_2) );
  AND2X1 gate2139 ( .A(N8387_1), .B(N8387_2), .Y(N8387) );
  AND2X1 gate2140 ( .A(N7020), .B(N4603), .Y(N8388) );
  AND2X1 gate2141_1 ( .A(N7036), .B(N7020), .Y(N8389_1) );
  AND2X1 gate2141 ( .A(N5981), .B(N8389_1), .Y(N8389) );
  AND2X1 gate2142 ( .A(N7020), .B(N4603), .Y(N8390) );
  AND2X1 gate2143_1 ( .A(N7036), .B(N7020), .Y(N8391_1) );
  AND2X1 gate2143 ( .A(N5981), .B(N8391_1), .Y(N8391) );
  AND2X1 gate2144 ( .A(N7036), .B(N5981), .Y(N8392) );
  AND2X1 gate2145 ( .A(N7049), .B(N6988), .Y(N8393) );
  AND2X1 gate2146 ( .A(N7057), .B(N7063), .Y(N8394) );
  AND2X1 gate2147 ( .A(N7057), .B(N7826), .Y(N8404) );
  AND2X1 gate2148_1 ( .A(N7098), .B(N7077), .Y(N8405_1) );
  AND2X1 gate2148_2 ( .A(N7073), .B(N7068), .Y(N8405_2) );
  AND2X1 gate2148 ( .A(N8405_1), .B(N8405_2), .Y(N8405) );
  AND2X1 gate2149 ( .A(N7068), .B(N4632), .Y(N8409) );
  AND2X1 gate2150_1 ( .A(N7073), .B(N7068), .Y(N8410_1) );
  AND2X1 gate2150 ( .A(N4634), .B(N8410_1), .Y(N8410) );
  AND2X1 gate2151_1 ( .A(N7077), .B(N7068), .Y(N8411_1) );
  AND2X1 gate2151_2 ( .A(N4635), .B(N7073), .Y(N8411_2) );
  AND2X1 gate2151 ( .A(N8411_1), .B(N8411_2), .Y(N8411) );
  AND2X1 gate2152_1 ( .A(N7099), .B(N7095), .Y(N8412_1) );
  AND2X1 gate2152_2 ( .A(N7091), .B(N7086), .Y(N8412_2) );
  AND2X1 gate2152_3 ( .A(N7080), .B(N8412_1), .Y(N8412_3) );
  AND2X1 gate2152 ( .A(N8412_2), .B(N8412_3), .Y(N8412) );
  AND2X1 gate2153 ( .A(N7080), .B(N4638), .Y(N8415) );
  AND2X1 gate2154_1 ( .A(N7086), .B(N7080), .Y(N8416_1) );
  AND2X1 gate2154 ( .A(N4639), .B(N8416_1), .Y(N8416) );
  AND2X1 gate2155_1 ( .A(N7091), .B(N7080), .Y(N8417_1) );
  AND2X1 gate2155_2 ( .A(N4640), .B(N7086), .Y(N8417_2) );
  AND2X1 gate2155 ( .A(N8417_1), .B(N8417_2), .Y(N8417) );
  AND2X1 gate2156_1 ( .A(N7095), .B(N7091), .Y(N8418_1) );
  AND2X1 gate2156_2 ( .A(N7080), .B(N4641), .Y(N8418_2) );
  AND2X1 gate2156_3 ( .A(N7086), .B(N8418_1), .Y(N8418_3) );
  AND2X1 gate2156 ( .A(N8418_2), .B(N8418_3), .Y(N8418) );
  AND2X1 gate2157 ( .A(N3375), .B(N7100), .Y(N8421) );
  AND2X1 gate2158_1 ( .A(N7114), .B(N7136), .Y(N8430_1) );
  AND2X1 gate2158_2 ( .A(N7125), .B(N7107), .Y(N8430_2) );
  AND2X1 gate2158 ( .A(N8430_1), .B(N8430_2), .Y(N8430) );
  AND2X1 gate2159 ( .A(N7107), .B(N4657), .Y(N8433) );
  AND2X1 gate2160_1 ( .A(N7114), .B(N7107), .Y(N8434_1) );
  AND2X1 gate2160 ( .A(N4661), .B(N8434_1), .Y(N8434) );
  AND2X1 gate2161_1 ( .A(N7125), .B(N7107), .Y(N8435_1) );
  AND2X1 gate2161_2 ( .A(N4667), .B(N7114), .Y(N8435_2) );
  AND2X1 gate2161 ( .A(N8435_1), .B(N8435_2), .Y(N8435) );
  AND2X1 gate2162 ( .A(N7114), .B(N4661), .Y(N8436) );
  AND2X1 gate2163_1 ( .A(N7125), .B(N4667), .Y(N8437_1) );
  AND2X1 gate2163 ( .A(N7114), .B(N8437_1), .Y(N8437) );
  AND2X1 gate2164_1 ( .A(N7136), .B(N7125), .Y(N8438_1) );
  AND2X1 gate2164 ( .A(N7114), .B(N8438_1), .Y(N8438) );
  AND2X1 gate2165 ( .A(N7114), .B(N4661), .Y(N8439) );
  AND2X1 gate2166_1 ( .A(N4667), .B(N7125), .Y(N8440_1) );
  AND2X1 gate2166 ( .A(N7114), .B(N8440_1), .Y(N8440) );
  AND2X1 gate2167 ( .A(N7125), .B(N4667), .Y(N8441) );
  AND2X1 gate2168 ( .A(N7136), .B(N7125), .Y(N8442) );
  AND2X1 gate2169 ( .A(N7125), .B(N4667), .Y(N8443) );
  AND2X1 gate2170_1 ( .A(N7149), .B(N7180), .Y(N8444_1) );
  AND2X1 gate2170_2 ( .A(N7159), .B(N7142), .Y(N8444_2) );
  AND2X1 gate2170_3 ( .A(N7170), .B(N8444_1), .Y(N8444_3) );
  AND2X1 gate2170 ( .A(N8444_2), .B(N8444_3), .Y(N8444) );
  AND2X1 gate2171 ( .A(N7142), .B(N4675), .Y(N8447) );
  AND2X1 gate2172_1 ( .A(N7149), .B(N7142), .Y(N8448_1) );
  AND2X1 gate2172 ( .A(N4678), .B(N8448_1), .Y(N8448) );
  AND2X1 gate2173_1 ( .A(N7159), .B(N7142), .Y(N8449_1) );
  AND2X1 gate2173_2 ( .A(N4682), .B(N7149), .Y(N8449_2) );
  AND2X1 gate2173 ( .A(N8449_1), .B(N8449_2), .Y(N8449) );
  AND2X1 gate2174_1 ( .A(N7170), .B(N7159), .Y(N8450_1) );
  AND2X1 gate2174_2 ( .A(N7142), .B(N4687), .Y(N8450_2) );
  AND2X1 gate2174_3 ( .A(N7149), .B(N8450_1), .Y(N8450_3) );
  AND2X1 gate2174 ( .A(N8450_2), .B(N8450_3), .Y(N8450) );
  AND2X1 gate2175 ( .A(N7149), .B(N4678), .Y(N8451) );
  AND2X1 gate2176_1 ( .A(N7159), .B(N4682), .Y(N8452_1) );
  AND2X1 gate2176 ( .A(N7149), .B(N8452_1), .Y(N8452) );
  AND2X1 gate2177_1 ( .A(N7170), .B(N7159), .Y(N8453_1) );
  AND2X1 gate2177_2 ( .A(N4687), .B(N7149), .Y(N8453_2) );
  AND2X1 gate2177 ( .A(N8453_1), .B(N8453_2), .Y(N8453) );
  AND2X1 gate2178 ( .A(N4682), .B(N7159), .Y(N8454) );
  AND2X1 gate2179_1 ( .A(N7170), .B(N7159), .Y(N8455_1) );
  AND2X1 gate2179 ( .A(N4687), .B(N8455_1), .Y(N8455) );
  AND2X1 gate2180 ( .A(N7170), .B(N4687), .Y(N8456) );
  INVX1 gate2181 ( .A(N7194), .Y(N8457) );
  INVX1 gate2182 ( .A(N7198), .Y(N8460) );
  INVX1 gate2183 ( .A(N7205), .Y(N8463) );
  INVX1 gate2184 ( .A(N7209), .Y(N8466) );
  INVX1 gate2185 ( .A(N7216), .Y(N8469) );
  INVX1 gate2186 ( .A(N7219), .Y(N8470) );
  BUFX2 gate2187 ( .A(N7202), .Y(N8471) );
  BUFX2 gate2188 ( .A(N7202), .Y(N8474) );
  BUFX2 gate2189 ( .A(N7213), .Y(N8477) );
  BUFX2 gate2190 ( .A(N7213), .Y(N8480) );
  AND2X1 gate2191_1 ( .A(N6083), .B(N6079), .Y(N8483_1) );
  AND2X1 gate2191 ( .A(N7216), .B(N8483_1), .Y(N8483) );
  AND2X1 gate2192_1 ( .A(N7191), .B(N7188), .Y(N8484_1) );
  AND2X1 gate2192 ( .A(N7219), .B(N8484_1), .Y(N8484) );
  AND2X1 gate2193_1 ( .A(N7301), .B(N7240), .Y(N8485_1) );
  AND2X1 gate2193_2 ( .A(N7229), .B(N7222), .Y(N8485_2) );
  AND2X1 gate2193 ( .A(N8485_1), .B(N8485_2), .Y(N8485) );
  AND2X1 gate2194 ( .A(N7222), .B(N4702), .Y(N8488) );
  AND2X1 gate2195_1 ( .A(N7229), .B(N7222), .Y(N8489_1) );
  AND2X1 gate2195 ( .A(N4706), .B(N8489_1), .Y(N8489) );
  AND2X1 gate2196_1 ( .A(N7240), .B(N7222), .Y(N8490_1) );
  AND2X1 gate2196_2 ( .A(N4711), .B(N7229), .Y(N8490_2) );
  AND2X1 gate2196 ( .A(N8490_1), .B(N8490_2), .Y(N8490) );
  AND2X1 gate2197 ( .A(N7229), .B(N4706), .Y(N8491) );
  AND2X1 gate2198_1 ( .A(N7240), .B(N4711), .Y(N8492_1) );
  AND2X1 gate2198 ( .A(N7229), .B(N8492_1), .Y(N8492) );
  AND2X1 gate2199_1 ( .A(N7301), .B(N7240), .Y(N8493_1) );
  AND2X1 gate2199 ( .A(N7229), .B(N8493_1), .Y(N8493) );
  AND2X1 gate2200 ( .A(N7229), .B(N4706), .Y(N8494) );
  AND2X1 gate2201_1 ( .A(N7240), .B(N4711), .Y(N8495_1) );
  AND2X1 gate2201 ( .A(N7229), .B(N8495_1), .Y(N8495) );
  AND2X1 gate2202 ( .A(N7240), .B(N4711), .Y(N8496) );
  AND2X1 gate2203_1 ( .A(N7307), .B(N7288), .Y(N8497_1) );
  AND2X1 gate2203_2 ( .A(N7272), .B(N7258), .Y(N8497_2) );
  AND2X1 gate2203_3 ( .A(N7250), .B(N8497_1), .Y(N8497_3) );
  AND2X1 gate2203 ( .A(N8497_2), .B(N8497_3), .Y(N8497) );
  AND2X1 gate2204 ( .A(N7250), .B(N4718), .Y(N8500) );
  AND2X1 gate2205_1 ( .A(N7258), .B(N7250), .Y(N8501_1) );
  AND2X1 gate2205 ( .A(N4722), .B(N8501_1), .Y(N8501) );
  AND2X1 gate2206_1 ( .A(N7272), .B(N7250), .Y(N8502_1) );
  AND2X1 gate2206_2 ( .A(N4728), .B(N7258), .Y(N8502_2) );
  AND2X1 gate2206 ( .A(N8502_1), .B(N8502_2), .Y(N8502) );
  AND2X1 gate2207_1 ( .A(N7288), .B(N7272), .Y(N8503_1) );
  AND2X1 gate2207_2 ( .A(N7250), .B(N4735), .Y(N8503_2) );
  AND2X1 gate2207_3 ( .A(N7258), .B(N8503_1), .Y(N8503_3) );
  AND2X1 gate2207 ( .A(N8503_2), .B(N8503_3), .Y(N8503) );
  AND2X1 gate2208 ( .A(N7258), .B(N4722), .Y(N8504) );
  AND2X1 gate2209_1 ( .A(N7272), .B(N4728), .Y(N8505_1) );
  AND2X1 gate2209 ( .A(N7258), .B(N8505_1), .Y(N8505) );
  AND2X1 gate2210_1 ( .A(N7288), .B(N7272), .Y(N8506_1) );
  AND2X1 gate2210_2 ( .A(N4735), .B(N7258), .Y(N8506_2) );
  AND2X1 gate2210 ( .A(N8506_1), .B(N8506_2), .Y(N8506) );
  AND2X1 gate2211_1 ( .A(N7307), .B(N7272), .Y(N8507_1) );
  AND2X1 gate2211_2 ( .A(N7258), .B(N7288), .Y(N8507_2) );
  AND2X1 gate2211 ( .A(N8507_1), .B(N8507_2), .Y(N8507) );
  AND2X1 gate2212 ( .A(N7258), .B(N4722), .Y(N8508) );
  AND2X1 gate2213_1 ( .A(N7272), .B(N4728), .Y(N8509_1) );
  AND2X1 gate2213 ( .A(N7258), .B(N8509_1), .Y(N8509) );
  AND2X1 gate2214_1 ( .A(N7288), .B(N7272), .Y(N8510_1) );
  AND2X1 gate2214_2 ( .A(N4735), .B(N7258), .Y(N8510_2) );
  AND2X1 gate2214 ( .A(N8510_1), .B(N8510_2), .Y(N8510) );
  AND2X1 gate2215 ( .A(N7272), .B(N4728), .Y(N8511) );
  AND2X1 gate2216_1 ( .A(N7288), .B(N7272), .Y(N8512_1) );
  AND2X1 gate2216 ( .A(N4735), .B(N8512_1), .Y(N8512) );
  AND2X1 gate2217_1 ( .A(N7307), .B(N7272), .Y(N8513_1) );
  AND2X1 gate2217 ( .A(N7288), .B(N8513_1), .Y(N8513) );
  AND2X1 gate2218 ( .A(N7272), .B(N4728), .Y(N8514) );
  AND2X1 gate2219_1 ( .A(N7288), .B(N7272), .Y(N8515_1) );
  AND2X1 gate2219 ( .A(N4735), .B(N8515_1), .Y(N8515) );
  AND2X1 gate2220 ( .A(N7288), .B(N4735), .Y(N8516) );
  AND2X1 gate2221 ( .A(N7301), .B(N7240), .Y(N8517) );
  AND2X1 gate2222 ( .A(N7307), .B(N7288), .Y(N8518) );
  INVX1 gate2223 ( .A(N7314), .Y(N8519) );
  INVX1 gate2224 ( .A(N7318), .Y(N8522) );
  BUFX2 gate2225 ( .A(N7322), .Y(N8525) );
  BUFX2 gate2226 ( .A(N7322), .Y(N8528) );
  BUFX2 gate2227 ( .A(N7331), .Y(N8531) );
  BUFX2 gate2228 ( .A(N7331), .Y(N8534) );
  INVX1 gate2229 ( .A(N7340), .Y(N8537) );
  INVX1 gate2230 ( .A(N7343), .Y(N8538) );
  AND2X1 gate2231_1 ( .A(N6141), .B(N6137), .Y(N8539_1) );
  AND2X1 gate2231 ( .A(N7340), .B(N8539_1), .Y(N8539) );
  AND2X1 gate2232_1 ( .A(N7337), .B(N7334), .Y(N8540_1) );
  AND2X1 gate2232 ( .A(N7343), .B(N8540_1), .Y(N8540) );
  AND2X1 gate2233_1 ( .A(N7376), .B(N7355), .Y(N8541_1) );
  AND2X1 gate2233_2 ( .A(N7351), .B(N7346), .Y(N8541_2) );
  AND2X1 gate2233 ( .A(N8541_1), .B(N8541_2), .Y(N8541) );
  AND2X1 gate2234 ( .A(N7346), .B(N4757), .Y(N8545) );
  AND2X1 gate2235_1 ( .A(N7351), .B(N7346), .Y(N8546_1) );
  AND2X1 gate2235 ( .A(N4758), .B(N8546_1), .Y(N8546) );
  AND2X1 gate2236_1 ( .A(N7355), .B(N7346), .Y(N8547_1) );
  AND2X1 gate2236_2 ( .A(N4759), .B(N7351), .Y(N8547_2) );
  AND2X1 gate2236 ( .A(N8547_1), .B(N8547_2), .Y(N8547) );
  AND2X1 gate2237_1 ( .A(N7377), .B(N7373), .Y(N8548_1) );
  AND2X1 gate2237_2 ( .A(N7369), .B(N7364), .Y(N8548_2) );
  AND2X1 gate2237_3 ( .A(N7358), .B(N8548_1), .Y(N8548_3) );
  AND2X1 gate2237 ( .A(N8548_2), .B(N8548_3), .Y(N8548) );
  AND2X1 gate2238 ( .A(N7358), .B(N4762), .Y(N8551) );
  AND2X1 gate2239_1 ( .A(N7364), .B(N7358), .Y(N8552_1) );
  AND2X1 gate2239 ( .A(N4764), .B(N8552_1), .Y(N8552) );
  AND2X1 gate2240_1 ( .A(N7369), .B(N7358), .Y(N8553_1) );
  AND2X1 gate2240_2 ( .A(N4766), .B(N7364), .Y(N8553_2) );
  AND2X1 gate2240 ( .A(N8553_1), .B(N8553_2), .Y(N8553) );
  AND2X1 gate2241_1 ( .A(N7373), .B(N7369), .Y(N8554_1) );
  AND2X1 gate2241_2 ( .A(N7358), .B(N4767), .Y(N8554_2) );
  AND2X1 gate2241_3 ( .A(N7364), .B(N8554_1), .Y(N8554_3) );
  AND2X1 gate2241 ( .A(N8554_2), .B(N8554_3), .Y(N8554) );
  INVX1 gate2242 ( .A(N7387), .Y(N8555) );
  INVX1 gate2243 ( .A(N7394), .Y(N8558) );
  INVX1 gate2244 ( .A(N7398), .Y(N8561) );
  INVX1 gate2245 ( .A(N7405), .Y(N8564) );
  INVX1 gate2246 ( .A(N7408), .Y(N8565) );
  BUFX2 gate2247 ( .A(N7391), .Y(N8566) );
  BUFX2 gate2248 ( .A(N7391), .Y(N8569) );
  BUFX2 gate2249 ( .A(N7402), .Y(N8572) );
  BUFX2 gate2250 ( .A(N7402), .Y(N8575) );
  AND2X1 gate2251_1 ( .A(N6170), .B(N6166), .Y(N8578_1) );
  AND2X1 gate2251 ( .A(N7405), .B(N8578_1), .Y(N8578) );
  AND2X1 gate2252_1 ( .A(N7381), .B(N7378), .Y(N8579_1) );
  AND2X1 gate2252 ( .A(N7408), .B(N8579_1), .Y(N8579) );
  BUFX2 gate2253 ( .A(N7180), .Y(N8580) );
  BUFX2 gate2254 ( .A(N7142), .Y(N8583) );
  BUFX2 gate2255 ( .A(N7149), .Y(N8586) );
  BUFX2 gate2256 ( .A(N7159), .Y(N8589) );
  BUFX2 gate2257 ( .A(N7170), .Y(N8592) );
  BUFX2 gate2258 ( .A(N6929), .Y(N8595) );
  BUFX2 gate2259 ( .A(N6936), .Y(N8598) );
  BUFX2 gate2260 ( .A(N6946), .Y(N8601) );
  BUFX2 gate2261 ( .A(N6957), .Y(N8604) );
  INVX1 gate2262 ( .A(N7441), .Y(N8607) );
  NAND2X1 gate2263 ( .A(N7441), .B(N5469), .Y(N8608) );
  INVX1 gate2264 ( .A(N7444), .Y(N8609) );
  NAND2X1 gate2265 ( .A(N7444), .B(N4793), .Y(N8610) );
  INVX1 gate2266 ( .A(N7447), .Y(N8615) );
  INVX1 gate2267 ( .A(N7450), .Y(N8616) );
  INVX1 gate2268 ( .A(N7453), .Y(N8617) );
  INVX1 gate2269 ( .A(N7456), .Y(N8618) );
  INVX1 gate2270 ( .A(N7474), .Y(N8619) );
  INVX1 gate2271 ( .A(N7465), .Y(N8624) );
  INVX1 gate2272 ( .A(N7468), .Y(N8625) );
  INVX1 gate2273 ( .A(N7471), .Y(N8626) );
  NAND2X1 gate2274 ( .A(N8144), .B(N8145), .Y(N8627) );
  INVX1 gate2275 ( .A(N7479), .Y(N8632) );
  INVX1 gate2276 ( .A(N7482), .Y(N8633) );
  INVX1 gate2277 ( .A(N7485), .Y(N8634) );
  INVX1 gate2278 ( .A(N7491), .Y(N8637) );
  INVX1 gate2279 ( .A(N7494), .Y(N8638) );
  INVX1 gate2280 ( .A(N7497), .Y(N8639) );
  INVX1 gate2281 ( .A(N7503), .Y(N8644) );
  INVX1 gate2282 ( .A(N7506), .Y(N8645) );
  INVX1 gate2283 ( .A(N7509), .Y(N8646) );
  INVX1 gate2284 ( .A(N7512), .Y(N8647) );
  INVX1 gate2285 ( .A(N7530), .Y(N8648) );
  INVX1 gate2286 ( .A(N7521), .Y(N8653) );
  INVX1 gate2287 ( .A(N7524), .Y(N8654) );
  INVX1 gate2288 ( .A(N7527), .Y(N8655) );
  BUFX2 gate2289 ( .A(N6894), .Y(N8660) );
  BUFX2 gate2290 ( .A(N6894), .Y(N8663) );
  BUFX2 gate2291 ( .A(N6901), .Y(N8666) );
  BUFX2 gate2292 ( .A(N6901), .Y(N8669) );
  BUFX2 gate2293 ( .A(N6912), .Y(N8672) );
  BUFX2 gate2294 ( .A(N6912), .Y(N8675) );
  BUFX2 gate2295 ( .A(N7049), .Y(N8678) );
  BUFX2 gate2296 ( .A(N6988), .Y(N8681) );
  BUFX2 gate2297 ( .A(N6970), .Y(N8684) );
  BUFX2 gate2298 ( .A(N6977), .Y(N8687) );
  BUFX2 gate2299 ( .A(N7049), .Y(N8690) );
  BUFX2 gate2300 ( .A(N6988), .Y(N8693) );
  BUFX2 gate2301 ( .A(N6970), .Y(N8696) );
  BUFX2 gate2302 ( .A(N6977), .Y(N8699) );
  BUFX2 gate2303 ( .A(N7036), .Y(N8702) );
  BUFX2 gate2304 ( .A(N6998), .Y(N8705) );
  BUFX2 gate2305 ( .A(N7020), .Y(N8708) );
  BUFX2 gate2306 ( .A(N7006), .Y(N8711) );
  BUFX2 gate2307 ( .A(N7006), .Y(N8714) );
  INVX1 gate2308 ( .A(N7553), .Y(N8717) );
  BUFX2 gate2309 ( .A(N7036), .Y(N8718) );
  BUFX2 gate2310 ( .A(N6998), .Y(N8721) );
  BUFX2 gate2311 ( .A(N7020), .Y(N8724) );
  NAND2X1 gate2312 ( .A(N8216), .B(N8217), .Y(N8727) );
  NAND2X1 gate2313 ( .A(N8218), .B(N8219), .Y(N8730) );
  INVX1 gate2314 ( .A(N7574), .Y(N8733) );
  INVX1 gate2315 ( .A(N7577), .Y(N8734) );
  BUFX2 gate2316 ( .A(N7107), .Y(N8735) );
  BUFX2 gate2317 ( .A(N7107), .Y(N8738) );
  BUFX2 gate2318 ( .A(N7114), .Y(N8741) );
  BUFX2 gate2319 ( .A(N7114), .Y(N8744) );
  BUFX2 gate2320 ( .A(N7125), .Y(N8747) );
  BUFX2 gate2321 ( .A(N7125), .Y(N8750) );
  INVX1 gate2322 ( .A(N7560), .Y(N8753) );
  INVX1 gate2323 ( .A(N7563), .Y(N8754) );
  INVX1 gate2324 ( .A(N7566), .Y(N8755) );
  INVX1 gate2325 ( .A(N7569), .Y(N8756) );
  BUFX2 gate2326 ( .A(N7301), .Y(N8757) );
  BUFX2 gate2327 ( .A(N7240), .Y(N8760) );
  BUFX2 gate2328 ( .A(N7222), .Y(N8763) );
  BUFX2 gate2329 ( .A(N7229), .Y(N8766) );
  BUFX2 gate2330 ( .A(N7301), .Y(N8769) );
  BUFX2 gate2331 ( .A(N7240), .Y(N8772) );
  BUFX2 gate2332 ( .A(N7222), .Y(N8775) );
  BUFX2 gate2333 ( .A(N7229), .Y(N8778) );
  BUFX2 gate2334 ( .A(N7307), .Y(N8781) );
  BUFX2 gate2335 ( .A(N7288), .Y(N8784) );
  BUFX2 gate2336 ( .A(N7250), .Y(N8787) );
  BUFX2 gate2337 ( .A(N7272), .Y(N8790) );
  BUFX2 gate2338 ( .A(N7258), .Y(N8793) );
  BUFX2 gate2339 ( .A(N7258), .Y(N8796) );
  BUFX2 gate2340 ( .A(N7307), .Y(N8799) );
  BUFX2 gate2341 ( .A(N7288), .Y(N8802) );
  BUFX2 gate2342 ( .A(N7250), .Y(N8805) );
  BUFX2 gate2343 ( .A(N7272), .Y(N8808) );
  NAND2X1 gate2344 ( .A(N8232), .B(N8233), .Y(N8811) );
  INVX1 gate2345 ( .A(N7588), .Y(N8814) );
  INVX1 gate2346 ( .A(N7591), .Y(N8815) );
  INVX1 gate2347 ( .A(N7582), .Y(N8816) );
  INVX1 gate2348 ( .A(N7585), .Y(N8817) );
  AND2X1 gate2349 ( .A(N7620), .B(N3155), .Y(N8818) );
  AND2X1 gate2350 ( .A(N3122), .B(N7609), .Y(N8840) );
  INVX1 gate2351 ( .A(N7609), .Y(N8857) );
  AND2X1 gate2352_1 ( .A(N6797), .B(N5740), .Y(N8861_1) );
  AND2X1 gate2352 ( .A(N8274), .B(N8861_1), .Y(N8861) );
  AND2X1 gate2353_1 ( .A(N5736), .B(N6800), .Y(N8862_1) );
  AND2X1 gate2353 ( .A(N8275), .B(N8862_1), .Y(N8862) );
  AND2X1 gate2354_1 ( .A(N6803), .B(N5751), .Y(N8863_1) );
  AND2X1 gate2354 ( .A(N8276), .B(N8863_1), .Y(N8863) );
  AND2X1 gate2355_1 ( .A(N5747), .B(N6806), .Y(N8864_1) );
  AND2X1 gate2355 ( .A(N8277), .B(N8864_1), .Y(N8864) );
  AND2X1 gate2356_1 ( .A(N6809), .B(N5762), .Y(N8865_1) );
  AND2X1 gate2356 ( .A(N8278), .B(N8865_1), .Y(N8865) );
  AND2X1 gate2357_1 ( .A(N5758), .B(N6812), .Y(N8866_1) );
  AND2X1 gate2357 ( .A(N8279), .B(N8866_1), .Y(N8866) );
  INVX1 gate2358 ( .A(N7655), .Y(N8871) );
  AND2X1 gate2359 ( .A(N6833), .B(N7655), .Y(N8874) );
  AND2X1 gate2360 ( .A(N7671), .B(N6867), .Y(N8878) );
  INVX1 gate2361 ( .A(N8196), .Y(N8879) );
  NAND2X1 gate2362 ( .A(N8196), .B(N8315), .Y(N8880) );
  INVX1 gate2363 ( .A(N8200), .Y(N8881) );
  NAND2X1 gate2364 ( .A(N8200), .B(N8317), .Y(N8882) );
  INVX1 gate2365 ( .A(N8204), .Y(N8883) );
  NAND2X1 gate2366 ( .A(N8204), .B(N8319), .Y(N8884) );
  INVX1 gate2367 ( .A(N8208), .Y(N8885) );
  NAND2X1 gate2368 ( .A(N8208), .B(N8321), .Y(N8886) );
  NAND2X1 gate2369 ( .A(N3658), .B(N8323), .Y(N8887) );
  NAND2X1 gate2370 ( .A(N4817), .B(N8325), .Y(N8888) );
  OR2X1 gate2371_1 ( .A(N4544), .B(N8337), .Y(N8898_1) );
  OR2X1 gate2371_2 ( .A(N8338), .B(N8339), .Y(N8898_2) );
  OR2X1 gate2371 ( .A(N8898_1), .B(N8898_2), .Y(N8898) );
  OR2X1 gate2372_1 ( .A(N4562), .B(N8348), .Y(N8902_1) );
  OR2X1 gate2372_2 ( .A(N8349), .B(N8350), .Y(N8902_2) );
  OR2X1 gate2372_3 ( .A(N8351), .B(N8902_1), .Y(N8902_3) );
  OR2X1 gate2372 ( .A(N8902_2), .B(N8902_3), .Y(N8902) );
  OR2X1 gate2373_1 ( .A(N4576), .B(N8369), .Y(N8920_1) );
  OR2X1 gate2373_2 ( .A(N8370), .B(N8371), .Y(N8920_2) );
  OR2X1 gate2373 ( .A(N8920_1), .B(N8920_2), .Y(N8920) );
  OR2X1 gate2374 ( .A(N4581), .B(N8377), .Y(N8924) );
  OR2X1 gate2375_1 ( .A(N4592), .B(N8378), .Y(N8927_1) );
  OR2X1 gate2375_2 ( .A(N8379), .B(N8380), .Y(N8927_2) );
  OR2X1 gate2375_3 ( .A(N8381), .B(N8927_1), .Y(N8927_3) );
  OR2X1 gate2375 ( .A(N8927_2), .B(N8927_3), .Y(N8927) );
  OR2X1 gate2376 ( .A(N4603), .B(N8392), .Y(N8931) );
  OR2X1 gate2377 ( .A(N7825), .B(N8404), .Y(N8943) );
  OR2X1 gate2378_1 ( .A(N4630), .B(N8409), .Y(N8950_1) );
  OR2X1 gate2378_2 ( .A(N8410), .B(N8411), .Y(N8950_2) );
  OR2X1 gate2378 ( .A(N8950_1), .B(N8950_2), .Y(N8950) );
  OR2X1 gate2379_1 ( .A(N4637), .B(N8415), .Y(N8956_1) );
  OR2X1 gate2379_2 ( .A(N8416), .B(N8417), .Y(N8956_2) );
  OR2X1 gate2379_3 ( .A(N8418), .B(N8956_1), .Y(N8956_3) );
  OR2X1 gate2379 ( .A(N8956_2), .B(N8956_3), .Y(N8956) );
  INVX1 gate2380 ( .A(N7852), .Y(N8959) );
  AND2X1 gate2381 ( .A(N3375), .B(N7852), .Y(N8960) );
  OR2X1 gate2382_1 ( .A(N4656), .B(N8433), .Y(N8963_1) );
  OR2X1 gate2382_2 ( .A(N8434), .B(N8435), .Y(N8963_2) );
  OR2X1 gate2382 ( .A(N8963_1), .B(N8963_2), .Y(N8963) );
  OR2X1 gate2383_1 ( .A(N4674), .B(N8447), .Y(N8966_1) );
  OR2X1 gate2383_2 ( .A(N8448), .B(N8449), .Y(N8966_2) );
  OR2X1 gate2383_3 ( .A(N8450), .B(N8966_1), .Y(N8966_3) );
  OR2X1 gate2383 ( .A(N8966_2), .B(N8966_3), .Y(N8966) );
  AND2X1 gate2384_1 ( .A(N7188), .B(N6083), .Y(N8991_1) );
  AND2X1 gate2384 ( .A(N8469), .B(N8991_1), .Y(N8991) );
  AND2X1 gate2385_1 ( .A(N6079), .B(N7191), .Y(N8992_1) );
  AND2X1 gate2385 ( .A(N8470), .B(N8992_1), .Y(N8992) );
  OR2X1 gate2386_1 ( .A(N4701), .B(N8488), .Y(N8995_1) );
  OR2X1 gate2386_2 ( .A(N8489), .B(N8490), .Y(N8995_2) );
  OR2X1 gate2386 ( .A(N8995_1), .B(N8995_2), .Y(N8995) );
  OR2X1 gate2387 ( .A(N4706), .B(N8496), .Y(N8996) );
  OR2X1 gate2388_1 ( .A(N4717), .B(N8500), .Y(N9001_1) );
  OR2X1 gate2388_2 ( .A(N8501), .B(N8502), .Y(N9001_2) );
  OR2X1 gate2388_3 ( .A(N8503), .B(N9001_1), .Y(N9001_3) );
  OR2X1 gate2388 ( .A(N9001_2), .B(N9001_3), .Y(N9001) );
  OR2X1 gate2389 ( .A(N4728), .B(N8516), .Y(N9005) );
  AND2X1 gate2390_1 ( .A(N7334), .B(N6141), .Y(N9024_1) );
  AND2X1 gate2390 ( .A(N8537), .B(N9024_1), .Y(N9024) );
  AND2X1 gate2391_1 ( .A(N6137), .B(N7337), .Y(N9025_1) );
  AND2X1 gate2391 ( .A(N8538), .B(N9025_1), .Y(N9025) );
  OR2X1 gate2392_1 ( .A(N4756), .B(N8545), .Y(N9029_1) );
  OR2X1 gate2392_2 ( .A(N8546), .B(N8547), .Y(N9029_2) );
  OR2X1 gate2392 ( .A(N9029_1), .B(N9029_2), .Y(N9029) );
  OR2X1 gate2393_1 ( .A(N4760), .B(N8551), .Y(N9035_1) );
  OR2X1 gate2393_2 ( .A(N8552), .B(N8553), .Y(N9035_2) );
  OR2X1 gate2393_3 ( .A(N8554), .B(N9035_1), .Y(N9035_3) );
  OR2X1 gate2393 ( .A(N9035_2), .B(N9035_3), .Y(N9035) );
  AND2X1 gate2394_1 ( .A(N7378), .B(N6170), .Y(N9053_1) );
  AND2X1 gate2394 ( .A(N8564), .B(N9053_1), .Y(N9053) );
  AND2X1 gate2395_1 ( .A(N6166), .B(N7381), .Y(N9054_1) );
  AND2X1 gate2395 ( .A(N8565), .B(N9054_1), .Y(N9054) );
  NAND2X1 gate2396 ( .A(N4303), .B(N8607), .Y(N9064) );
  NAND2X1 gate2397 ( .A(N3507), .B(N8609), .Y(N9065) );
  INVX1 gate2398 ( .A(N8114), .Y(N9066) );
  NAND2X1 gate2399 ( .A(N8114), .B(N4795), .Y(N9067) );
  OR2X1 gate2400 ( .A(N7613), .B(N6783), .Y(N9068) );
  INVX1 gate2401 ( .A(N8117), .Y(N9071) );
  INVX1 gate2402 ( .A(N8131), .Y(N9072) );
  NAND2X1 gate2403 ( .A(N8131), .B(N6195), .Y(N9073) );
  INVX1 gate2404 ( .A(N7613), .Y(N9074) );
  INVX1 gate2405 ( .A(N8134), .Y(N9077) );
  OR2X1 gate2406 ( .A(N7650), .B(N6865), .Y(N9079) );
  INVX1 gate2407 ( .A(N8146), .Y(N9082) );
  INVX1 gate2408 ( .A(N7650), .Y(N9083) );
  INVX1 gate2409 ( .A(N8156), .Y(N9086) );
  INVX1 gate2410 ( .A(N8166), .Y(N9087) );
  NAND2X1 gate2411 ( .A(N8166), .B(N4813), .Y(N9088) );
  OR2X1 gate2412 ( .A(N7659), .B(N6866), .Y(N9089) );
  INVX1 gate2413 ( .A(N8169), .Y(N9092) );
  INVX1 gate2414 ( .A(N8183), .Y(N9093) );
  NAND2X1 gate2415 ( .A(N8183), .B(N6203), .Y(N9094) );
  INVX1 gate2416 ( .A(N7659), .Y(N9095) );
  INVX1 gate2417 ( .A(N8186), .Y(N9098) );
  OR2X1 gate2418_1 ( .A(N4545), .B(N8340), .Y(N9099_1) );
  OR2X1 gate2418_2 ( .A(N8341), .B(N8342), .Y(N9099_2) );
  OR2X1 gate2418 ( .A(N9099_1), .B(N9099_2), .Y(N9099) );
  NOR3X1 gate2419 ( .A(N4545), .B(N8343), .C(N8344), .Y(N9103) );
  OR2X1 gate2420_1 ( .A(N4549), .B(N8345), .Y(N9107_1) );
  OR2X1 gate2420 ( .A(N8346), .B(N9107_1), .Y(N9107) );
  NOR2X1 gate2421 ( .A(N4549), .B(N8347), .Y(N9111) );
  OR2X1 gate2422_1 ( .A(N4577), .B(N8372), .Y(N9117_1) );
  OR2X1 gate2422_2 ( .A(N8373), .B(N8374), .Y(N9117_2) );
  OR2X1 gate2422 ( .A(N9117_1), .B(N9117_2), .Y(N9117) );
  NOR3X1 gate2423 ( .A(N4577), .B(N8375), .C(N8376), .Y(N9127) );
  NOR3X1 gate2424 ( .A(N4597), .B(N8390), .C(N8391), .Y(N9146) );
  NOR2X1 gate2425_1 ( .A(N4593), .B(N8385), .Y(N9149_1) );
  NOR2X1 gate2425_2 ( .A(N8386), .B(N8387), .Y(N9149_2) );
  NOR2X1 gate2425 ( .A(N9149_1), .B(N9149_2), .Y(N9149) );
  NAND2X1 gate2426 ( .A(N7577), .B(N8733), .Y(N9159) );
  NAND2X1 gate2427 ( .A(N7574), .B(N8734), .Y(N9160) );
  OR2X1 gate2428_1 ( .A(N4657), .B(N8436), .Y(N9161_1) );
  OR2X1 gate2428_2 ( .A(N8437), .B(N8438), .Y(N9161_2) );
  OR2X1 gate2428 ( .A(N9161_1), .B(N9161_2), .Y(N9161) );
  NOR3X1 gate2429 ( .A(N4657), .B(N8439), .C(N8440), .Y(N9165) );
  OR2X1 gate2430_1 ( .A(N4661), .B(N8441), .Y(N9169_1) );
  OR2X1 gate2430 ( .A(N8442), .B(N9169_1), .Y(N9169) );
  NOR2X1 gate2431 ( .A(N4661), .B(N8443), .Y(N9173) );
  NAND2X1 gate2432 ( .A(N7563), .B(N8753), .Y(N9179) );
  NAND2X1 gate2433 ( .A(N7560), .B(N8754), .Y(N9180) );
  NAND2X1 gate2434 ( .A(N7569), .B(N8755), .Y(N9181) );
  NAND2X1 gate2435 ( .A(N7566), .B(N8756), .Y(N9182) );
  OR2X1 gate2436_1 ( .A(N4702), .B(N8491), .Y(N9183_1) );
  OR2X1 gate2436_2 ( .A(N8492), .B(N8493), .Y(N9183_2) );
  OR2X1 gate2436 ( .A(N9183_1), .B(N9183_2), .Y(N9183) );
  NOR3X1 gate2437 ( .A(N4702), .B(N8494), .C(N8495), .Y(N9193) );
  OR2X1 gate2438_1 ( .A(N4722), .B(N8511), .Y(N9203_1) );
  OR2X1 gate2438_2 ( .A(N8512), .B(N8513), .Y(N9203_2) );
  OR2X1 gate2438 ( .A(N9203_1), .B(N9203_2), .Y(N9203) );
  OR2X1 gate2439_1 ( .A(N4718), .B(N8504), .Y(N9206_1) );
  OR2X1 gate2439_2 ( .A(N8505), .B(N8506), .Y(N9206_2) );
  OR2X1 gate2439_3 ( .A(N8507), .B(N9206_1), .Y(N9206_3) );
  OR2X1 gate2439 ( .A(N9206_2), .B(N9206_3), .Y(N9206) );
  NOR3X1 gate2440 ( .A(N4722), .B(N8514), .C(N8515), .Y(N9220) );
  NOR2X1 gate2441_1 ( .A(N4718), .B(N8508), .Y(N9223_1) );
  NOR2X1 gate2441_2 ( .A(N8509), .B(N8510), .Y(N9223_2) );
  NOR2X1 gate2441 ( .A(N9223_1), .B(N9223_2), .Y(N9223) );
  NAND2X1 gate2442 ( .A(N7591), .B(N8814), .Y(N9234) );
  NAND2X1 gate2443 ( .A(N7588), .B(N8815), .Y(N9235) );
  NAND2X1 gate2444 ( .A(N7585), .B(N8816), .Y(N9236) );
  NAND2X1 gate2445 ( .A(N7582), .B(N8817), .Y(N9237) );
  OR2X1 gate2446 ( .A(N3159), .B(N8818), .Y(N9238) );
  OR2X1 gate2447 ( .A(N3126), .B(N8840), .Y(N9242) );
  NAND2X1 gate2448 ( .A(N8324), .B(N8888), .Y(N9243) );
  INVX1 gate2449 ( .A(N8580), .Y(N9244) );
  INVX1 gate2450 ( .A(N8583), .Y(N9245) );
  INVX1 gate2451 ( .A(N8586), .Y(N9246) );
  INVX1 gate2452 ( .A(N8589), .Y(N9247) );
  INVX1 gate2453 ( .A(N8592), .Y(N9248) );
  INVX1 gate2454 ( .A(N8595), .Y(N9249) );
  INVX1 gate2455 ( .A(N8598), .Y(N9250) );
  INVX1 gate2456 ( .A(N8601), .Y(N9251) );
  INVX1 gate2457 ( .A(N8604), .Y(N9252) );
  NOR2X1 gate2458 ( .A(N8861), .B(N8280), .Y(N9256) );
  NOR2X1 gate2459 ( .A(N8862), .B(N8281), .Y(N9257) );
  NOR2X1 gate2460 ( .A(N8863), .B(N8282), .Y(N9258) );
  NOR2X1 gate2461 ( .A(N8864), .B(N8283), .Y(N9259) );
  NOR2X1 gate2462 ( .A(N8865), .B(N8284), .Y(N9260) );
  NOR2X1 gate2463 ( .A(N8866), .B(N8285), .Y(N9261) );
  INVX1 gate2464 ( .A(N8627), .Y(N9262) );
  OR2X1 gate2465 ( .A(N7649), .B(N8874), .Y(N9265) );
  OR2X1 gate2466 ( .A(N7668), .B(N8878), .Y(N9268) );
  NAND2X1 gate2467 ( .A(N7533), .B(N8879), .Y(N9271) );
  NAND2X1 gate2468 ( .A(N7536), .B(N8881), .Y(N9272) );
  NAND2X1 gate2469 ( .A(N7539), .B(N8883), .Y(N9273) );
  NAND2X1 gate2470 ( .A(N7542), .B(N8885), .Y(N9274) );
  NAND2X1 gate2471 ( .A(N8322), .B(N8887), .Y(N9275) );
  INVX1 gate2472 ( .A(N8333), .Y(N9276) );
  AND2X1 gate2473_1 ( .A(N6936), .B(N8326), .Y(N9280_1) );
  AND2X1 gate2473_2 ( .A(N6946), .B(N6929), .Y(N9280_2) );
  AND2X1 gate2473_3 ( .A(N6957), .B(N9280_1), .Y(N9280_3) );
  AND2X1 gate2473 ( .A(N9280_2), .B(N9280_3), .Y(N9280) );
  AND2X1 gate2474_1 ( .A(N367), .B(N8326), .Y(N9285_1) );
  AND2X1 gate2474_2 ( .A(N6946), .B(N6957), .Y(N9285_2) );
  AND2X1 gate2474_3 ( .A(N6936), .B(N9285_1), .Y(N9285_3) );
  AND2X1 gate2474 ( .A(N9285_2), .B(N9285_3), .Y(N9285) );
  AND2X1 gate2475_1 ( .A(N367), .B(N8326), .Y(N9286_1) );
  AND2X1 gate2475_2 ( .A(N6946), .B(N6957), .Y(N9286_2) );
  AND2X1 gate2475 ( .A(N9286_1), .B(N9286_2), .Y(N9286) );
  AND2X1 gate2476_1 ( .A(N367), .B(N8326), .Y(N9287_1) );
  AND2X1 gate2476 ( .A(N6957), .B(N9287_1), .Y(N9287) );
  AND2X1 gate2477 ( .A(N367), .B(N8326), .Y(N9288) );
  INVX1 gate2478 ( .A(N8660), .Y(N9290) );
  INVX1 gate2479 ( .A(N8663), .Y(N9292) );
  INVX1 gate2480 ( .A(N8666), .Y(N9294) );
  INVX1 gate2481 ( .A(N8669), .Y(N9296) );
  NAND2X1 gate2482 ( .A(N8672), .B(N5966), .Y(N9297) );
  INVX1 gate2483 ( .A(N8672), .Y(N9298) );
  NAND2X1 gate2484 ( .A(N8675), .B(N6969), .Y(N9299) );
  INVX1 gate2485 ( .A(N8675), .Y(N9300) );
  INVX1 gate2486 ( .A(N8365), .Y(N9301) );
  AND2X1 gate2487_1 ( .A(N8358), .B(N7036), .Y(N9307_1) );
  AND2X1 gate2487_2 ( .A(N7020), .B(N7006), .Y(N9307_2) );
  AND2X1 gate2487_3 ( .A(N6998), .B(N9307_1), .Y(N9307_3) );
  AND2X1 gate2487 ( .A(N9307_2), .B(N9307_3), .Y(N9307) );
  AND2X1 gate2488_1 ( .A(N8358), .B(N7020), .Y(N9314_1) );
  AND2X1 gate2488_2 ( .A(N7006), .B(N7036), .Y(N9314_2) );
  AND2X1 gate2488 ( .A(N9314_1), .B(N9314_2), .Y(N9314) );
  AND2X1 gate2489_1 ( .A(N8358), .B(N7020), .Y(N9315_1) );
  AND2X1 gate2489 ( .A(N7036), .B(N9315_1), .Y(N9315) );
  AND2X1 gate2490 ( .A(N8358), .B(N7036), .Y(N9318) );
  INVX1 gate2491 ( .A(N8687), .Y(N9319) );
  INVX1 gate2492 ( .A(N8699), .Y(N9320) );
  INVX1 gate2493 ( .A(N8711), .Y(N9321) );
  INVX1 gate2494 ( .A(N8714), .Y(N9322) );
  INVX1 gate2495 ( .A(N8727), .Y(N9323) );
  INVX1 gate2496 ( .A(N8730), .Y(N9324) );
  INVX1 gate2497 ( .A(N8405), .Y(N9326) );
  AND2X1 gate2498 ( .A(N8405), .B(N8412), .Y(N9332) );
  OR2X1 gate2499 ( .A(N4193), .B(N8960), .Y(N9339) );
  AND2X1 gate2500 ( .A(N8430), .B(N8444), .Y(N9344) );
  INVX1 gate2501 ( .A(N8735), .Y(N9352) );
  INVX1 gate2502 ( .A(N8738), .Y(N9354) );
  INVX1 gate2503 ( .A(N8741), .Y(N9356) );
  INVX1 gate2504 ( .A(N8744), .Y(N9358) );
  NAND2X1 gate2505 ( .A(N8747), .B(N6078), .Y(N9359) );
  INVX1 gate2506 ( .A(N8747), .Y(N9360) );
  NAND2X1 gate2507 ( .A(N8750), .B(N7187), .Y(N9361) );
  INVX1 gate2508 ( .A(N8750), .Y(N9362) );
  INVX1 gate2509 ( .A(N8471), .Y(N9363) );
  INVX1 gate2510 ( .A(N8474), .Y(N9364) );
  INVX1 gate2511 ( .A(N8477), .Y(N9365) );
  INVX1 gate2512 ( .A(N8480), .Y(N9366) );
  NOR2X1 gate2513 ( .A(N8991), .B(N8483), .Y(N9367) );
  NOR2X1 gate2514 ( .A(N8992), .B(N8484), .Y(N9368) );
  AND2X1 gate2515_1 ( .A(N7198), .B(N7194), .Y(N9369_1) );
  AND2X1 gate2515 ( .A(N8471), .B(N9369_1), .Y(N9369) );
  AND2X1 gate2516_1 ( .A(N8460), .B(N8457), .Y(N9370_1) );
  AND2X1 gate2516 ( .A(N8474), .B(N9370_1), .Y(N9370) );
  AND2X1 gate2517_1 ( .A(N7209), .B(N7205), .Y(N9371_1) );
  AND2X1 gate2517 ( .A(N8477), .B(N9371_1), .Y(N9371) );
  AND2X1 gate2518_1 ( .A(N8466), .B(N8463), .Y(N9372_1) );
  AND2X1 gate2518 ( .A(N8480), .B(N9372_1), .Y(N9372) );
  INVX1 gate2519 ( .A(N8497), .Y(N9375) );
  INVX1 gate2520 ( .A(N8766), .Y(N9381) );
  INVX1 gate2521 ( .A(N8778), .Y(N9382) );
  INVX1 gate2522 ( .A(N8793), .Y(N9383) );
  INVX1 gate2523 ( .A(N8796), .Y(N9384) );
  AND2X1 gate2524 ( .A(N8485), .B(N8497), .Y(N9385) );
  INVX1 gate2525 ( .A(N8525), .Y(N9392) );
  INVX1 gate2526 ( .A(N8528), .Y(N9393) );
  INVX1 gate2527 ( .A(N8531), .Y(N9394) );
  INVX1 gate2528 ( .A(N8534), .Y(N9395) );
  AND2X1 gate2529_1 ( .A(N7318), .B(N7314), .Y(N9396_1) );
  AND2X1 gate2529 ( .A(N8525), .B(N9396_1), .Y(N9396) );
  AND2X1 gate2530_1 ( .A(N8522), .B(N8519), .Y(N9397_1) );
  AND2X1 gate2530 ( .A(N8528), .B(N9397_1), .Y(N9397) );
  AND2X1 gate2531_1 ( .A(N6131), .B(N6127), .Y(N9398_1) );
  AND2X1 gate2531 ( .A(N8531), .B(N9398_1), .Y(N9398) );
  AND2X1 gate2532_1 ( .A(N7328), .B(N7325), .Y(N9399_1) );
  AND2X1 gate2532 ( .A(N8534), .B(N9399_1), .Y(N9399) );
  NOR2X1 gate2533 ( .A(N9024), .B(N8539), .Y(N9400) );
  NOR2X1 gate2534 ( .A(N9025), .B(N8540), .Y(N9401) );
  INVX1 gate2535 ( .A(N8541), .Y(N9402) );
  NAND2X1 gate2536 ( .A(N8548), .B(N89), .Y(N9407) );
  AND2X1 gate2537 ( .A(N8541), .B(N8548), .Y(N9408) );
  INVX1 gate2538 ( .A(N8811), .Y(N9412) );
  INVX1 gate2539 ( .A(N8566), .Y(N9413) );
  INVX1 gate2540 ( .A(N8569), .Y(N9414) );
  INVX1 gate2541 ( .A(N8572), .Y(N9415) );
  INVX1 gate2542 ( .A(N8575), .Y(N9416) );
  NOR2X1 gate2543 ( .A(N9053), .B(N8578), .Y(N9417) );
  NOR2X1 gate2544 ( .A(N9054), .B(N8579), .Y(N9418) );
  AND2X1 gate2545_1 ( .A(N7387), .B(N6177), .Y(N9419_1) );
  AND2X1 gate2545 ( .A(N8566), .B(N9419_1), .Y(N9419) );
  AND2X1 gate2546_1 ( .A(N8555), .B(N7384), .Y(N9420_1) );
  AND2X1 gate2546 ( .A(N8569), .B(N9420_1), .Y(N9420) );
  AND2X1 gate2547_1 ( .A(N7398), .B(N7394), .Y(N9421_1) );
  AND2X1 gate2547 ( .A(N8572), .B(N9421_1), .Y(N9421) );
  AND2X1 gate2548_1 ( .A(N8561), .B(N8558), .Y(N9422_1) );
  AND2X1 gate2548 ( .A(N8575), .B(N9422_1), .Y(N9422) );
  BUFX2 gate2549 ( .A(N8326), .Y(N9423) );
  NAND2X1 gate2550 ( .A(N9064), .B(N8608), .Y(N9426) );
  NAND2X1 gate2551 ( .A(N9065), .B(N8610), .Y(N9429) );
  NAND2X1 gate2552 ( .A(N3515), .B(N9066), .Y(N9432) );
  NAND2X1 gate2553 ( .A(N4796), .B(N9072), .Y(N9435) );
  NAND2X1 gate2554 ( .A(N3628), .B(N9087), .Y(N9442) );
  NAND2X1 gate2555 ( .A(N4814), .B(N9093), .Y(N9445) );
  INVX1 gate2556 ( .A(N8678), .Y(N9454) );
  INVX1 gate2557 ( .A(N8681), .Y(N9455) );
  INVX1 gate2558 ( .A(N8684), .Y(N9456) );
  INVX1 gate2559 ( .A(N8690), .Y(N9459) );
  INVX1 gate2560 ( .A(N8693), .Y(N9460) );
  INVX1 gate2561 ( .A(N8696), .Y(N9461) );
  BUFX2 gate2562 ( .A(N8358), .Y(N9462) );
  INVX1 gate2563 ( .A(N8702), .Y(N9465) );
  INVX1 gate2564 ( .A(N8705), .Y(N9466) );
  INVX1 gate2565 ( .A(N8708), .Y(N9467) );
  INVX1 gate2566 ( .A(N8724), .Y(N9468) );
  BUFX2 gate2567 ( .A(N8358), .Y(N9473) );
  INVX1 gate2568 ( .A(N8718), .Y(N9476) );
  INVX1 gate2569 ( .A(N8721), .Y(N9477) );
  NAND2X1 gate2570 ( .A(N9159), .B(N9160), .Y(N9478) );
  NAND2X1 gate2571 ( .A(N9179), .B(N9180), .Y(N9485) );
  NAND2X1 gate2572 ( .A(N9181), .B(N9182), .Y(N9488) );
  INVX1 gate2573 ( .A(N8757), .Y(N9493) );
  INVX1 gate2574 ( .A(N8760), .Y(N9494) );
  INVX1 gate2575 ( .A(N8763), .Y(N9495) );
  INVX1 gate2576 ( .A(N8769), .Y(N9498) );
  INVX1 gate2577 ( .A(N8772), .Y(N9499) );
  INVX1 gate2578 ( .A(N8775), .Y(N9500) );
  INVX1 gate2579 ( .A(N8781), .Y(N9505) );
  INVX1 gate2580 ( .A(N8784), .Y(N9506) );
  INVX1 gate2581 ( .A(N8787), .Y(N9507) );
  INVX1 gate2582 ( .A(N8790), .Y(N9508) );
  INVX1 gate2583 ( .A(N8808), .Y(N9509) );
  INVX1 gate2584 ( .A(N8799), .Y(N9514) );
  INVX1 gate2585 ( .A(N8802), .Y(N9515) );
  INVX1 gate2586 ( .A(N8805), .Y(N9516) );
  NAND2X1 gate2587 ( .A(N9234), .B(N9235), .Y(N9517) );
  NAND2X1 gate2588 ( .A(N9236), .B(N9237), .Y(N9520) );
  AND2X1 gate2589 ( .A(N8943), .B(N8421), .Y(N9526) );
  AND2X1 gate2590 ( .A(N8943), .B(N8421), .Y(N9531) );
  NAND2X1 gate2591 ( .A(N9271), .B(N8880), .Y(N9539) );
  NAND2X1 gate2592 ( .A(N9273), .B(N8884), .Y(N9540) );
  INVX1 gate2593 ( .A(N9275), .Y(N9541) );
  AND2X1 gate2594 ( .A(N8857), .B(N8254), .Y(N9543) );
  AND2X1 gate2595 ( .A(N8871), .B(N8288), .Y(N9551) );
  NAND2X1 gate2596 ( .A(N9272), .B(N8882), .Y(N9555) );
  NAND2X1 gate2597 ( .A(N9274), .B(N8886), .Y(N9556) );
  INVX1 gate2598 ( .A(N8898), .Y(N9557) );
  AND2X1 gate2599 ( .A(N8902), .B(N8333), .Y(N9560) );
  INVX1 gate2600 ( .A(N9099), .Y(N9561) );
  NAND2X1 gate2601 ( .A(N9099), .B(N9290), .Y(N9562) );
  INVX1 gate2602 ( .A(N9103), .Y(N9563) );
  NAND2X1 gate2603 ( .A(N9103), .B(N9292), .Y(N9564) );
  INVX1 gate2604 ( .A(N9107), .Y(N9565) );
  NAND2X1 gate2605 ( .A(N9107), .B(N9294), .Y(N9566) );
  INVX1 gate2606 ( .A(N9111), .Y(N9567) );
  NAND2X1 gate2607 ( .A(N9111), .B(N9296), .Y(N9568) );
  NAND2X1 gate2608 ( .A(N4844), .B(N9298), .Y(N9569) );
  NAND2X1 gate2609 ( .A(N6207), .B(N9300), .Y(N9570) );
  INVX1 gate2610 ( .A(N8920), .Y(N9571) );
  INVX1 gate2611 ( .A(N8927), .Y(N9575) );
  AND2X1 gate2612 ( .A(N8365), .B(N8927), .Y(N9579) );
  INVX1 gate2613 ( .A(N8950), .Y(N9581) );
  INVX1 gate2614 ( .A(N8956), .Y(N9582) );
  AND2X1 gate2615 ( .A(N8405), .B(N8956), .Y(N9585) );
  AND2X1 gate2616 ( .A(N8966), .B(N8430), .Y(N9591) );
  INVX1 gate2617 ( .A(N9161), .Y(N9592) );
  NAND2X1 gate2618 ( .A(N9161), .B(N9352), .Y(N9593) );
  INVX1 gate2619 ( .A(N9165), .Y(N9594) );
  NAND2X1 gate2620 ( .A(N9165), .B(N9354), .Y(N9595) );
  INVX1 gate2621 ( .A(N9169), .Y(N9596) );
  NAND2X1 gate2622 ( .A(N9169), .B(N9356), .Y(N9597) );
  INVX1 gate2623 ( .A(N9173), .Y(N9598) );
  NAND2X1 gate2624 ( .A(N9173), .B(N9358), .Y(N9599) );
  NAND2X1 gate2625 ( .A(N4940), .B(N9360), .Y(N9600) );
  NAND2X1 gate2626 ( .A(N6220), .B(N9362), .Y(N9601) );
  AND2X1 gate2627_1 ( .A(N8457), .B(N7198), .Y(N9602_1) );
  AND2X1 gate2627 ( .A(N9363), .B(N9602_1), .Y(N9602) );
  AND2X1 gate2628_1 ( .A(N7194), .B(N8460), .Y(N9603_1) );
  AND2X1 gate2628 ( .A(N9364), .B(N9603_1), .Y(N9603) );
  AND2X1 gate2629_1 ( .A(N8463), .B(N7209), .Y(N9604_1) );
  AND2X1 gate2629 ( .A(N9365), .B(N9604_1), .Y(N9604) );
  AND2X1 gate2630_1 ( .A(N7205), .B(N8466), .Y(N9605_1) );
  AND2X1 gate2630 ( .A(N9366), .B(N9605_1), .Y(N9605) );
  INVX1 gate2631 ( .A(N9001), .Y(N9608) );
  AND2X1 gate2632 ( .A(N8485), .B(N9001), .Y(N9611) );
  AND2X1 gate2633_1 ( .A(N8519), .B(N7318), .Y(N9612_1) );
  AND2X1 gate2633 ( .A(N9392), .B(N9612_1), .Y(N9612) );
  AND2X1 gate2634_1 ( .A(N7314), .B(N8522), .Y(N9613_1) );
  AND2X1 gate2634 ( .A(N9393), .B(N9613_1), .Y(N9613) );
  AND2X1 gate2635_1 ( .A(N7325), .B(N6131), .Y(N9614_1) );
  AND2X1 gate2635 ( .A(N9394), .B(N9614_1), .Y(N9614) );
  AND2X1 gate2636_1 ( .A(N6127), .B(N7328), .Y(N9615_1) );
  AND2X1 gate2636 ( .A(N9395), .B(N9615_1), .Y(N9615) );
  INVX1 gate2637 ( .A(N9029), .Y(N9616) );
  INVX1 gate2638 ( .A(N9035), .Y(N9617) );
  AND2X1 gate2639 ( .A(N8541), .B(N9035), .Y(N9618) );
  AND2X1 gate2640_1 ( .A(N7384), .B(N7387), .Y(N9621_1) );
  AND2X1 gate2640 ( .A(N9413), .B(N9621_1), .Y(N9621) );
  AND2X1 gate2641_1 ( .A(N6177), .B(N8555), .Y(N9622_1) );
  AND2X1 gate2641 ( .A(N9414), .B(N9622_1), .Y(N9622) );
  AND2X1 gate2642_1 ( .A(N8558), .B(N7398), .Y(N9623_1) );
  AND2X1 gate2642 ( .A(N9415), .B(N9623_1), .Y(N9623) );
  AND2X1 gate2643_1 ( .A(N7394), .B(N8561), .Y(N9624_1) );
  AND2X1 gate2643 ( .A(N9416), .B(N9624_1), .Y(N9624) );
  OR2X1 gate2644_1 ( .A(N4563), .B(N8352), .Y(N9626_1) );
  OR2X1 gate2644_2 ( .A(N8353), .B(N8354), .Y(N9626_2) );
  OR2X1 gate2644_3 ( .A(N9285), .B(N9626_1), .Y(N9626_3) );
  OR2X1 gate2644 ( .A(N9626_2), .B(N9626_3), .Y(N9626) );
  OR2X1 gate2645_1 ( .A(N4566), .B(N8355), .Y(N9629_1) );
  OR2X1 gate2645_2 ( .A(N8356), .B(N9286), .Y(N9629_2) );
  OR2X1 gate2645 ( .A(N9629_1), .B(N9629_2), .Y(N9629) );
  OR2X1 gate2646_1 ( .A(N4570), .B(N8357), .Y(N9632_1) );
  OR2X1 gate2646 ( .A(N9287), .B(N9632_1), .Y(N9632) );
  OR2X1 gate2647 ( .A(N5960), .B(N9288), .Y(N9635) );
  NAND2X1 gate2648 ( .A(N9067), .B(N9432), .Y(N9642) );
  INVX1 gate2649 ( .A(N9068), .Y(N9645) );
  NAND2X1 gate2650 ( .A(N9073), .B(N9435), .Y(N9646) );
  INVX1 gate2651 ( .A(N9074), .Y(N9649) );
  NAND2X1 gate2652 ( .A(N9257), .B(N9256), .Y(N9650) );
  NAND2X1 gate2653 ( .A(N9259), .B(N9258), .Y(N9653) );
  NAND2X1 gate2654 ( .A(N9261), .B(N9260), .Y(N9656) );
  INVX1 gate2655 ( .A(N9079), .Y(N9659) );
  NAND2X1 gate2656 ( .A(N9079), .B(N4809), .Y(N9660) );
  INVX1 gate2657 ( .A(N9083), .Y(N9661) );
  NAND2X1 gate2658 ( .A(N9083), .B(N6202), .Y(N9662) );
  NAND2X1 gate2659 ( .A(N9088), .B(N9442), .Y(N9663) );
  INVX1 gate2660 ( .A(N9089), .Y(N9666) );
  NAND2X1 gate2661 ( .A(N9094), .B(N9445), .Y(N9667) );
  INVX1 gate2662 ( .A(N9095), .Y(N9670) );
  OR2X1 gate2663 ( .A(N8924), .B(N8393), .Y(N9671) );
  INVX1 gate2664 ( .A(N9117), .Y(N9674) );
  INVX1 gate2665 ( .A(N8924), .Y(N9675) );
  INVX1 gate2666 ( .A(N9127), .Y(N9678) );
  OR2X1 gate2667_1 ( .A(N4597), .B(N8388), .Y(N9679_1) );
  OR2X1 gate2667_2 ( .A(N8389), .B(N9315), .Y(N9679_2) );
  OR2X1 gate2667 ( .A(N9679_1), .B(N9679_2), .Y(N9679) );
  OR2X1 gate2668 ( .A(N8931), .B(N9318), .Y(N9682) );
  OR2X1 gate2669_1 ( .A(N4593), .B(N8382), .Y(N9685_1) );
  OR2X1 gate2669_2 ( .A(N8383), .B(N8384), .Y(N9685_2) );
  OR2X1 gate2669_3 ( .A(N9314), .B(N9685_1), .Y(N9685_3) );
  OR2X1 gate2669 ( .A(N9685_2), .B(N9685_3), .Y(N9685) );
  INVX1 gate2670 ( .A(N9146), .Y(N9690) );
  NAND2X1 gate2671 ( .A(N9146), .B(N8717), .Y(N9691) );
  INVX1 gate2672 ( .A(N8931), .Y(N9692) );
  INVX1 gate2673 ( .A(N9149), .Y(N9695) );
  NAND2X1 gate2674 ( .A(N9401), .B(N9400), .Y(N9698) );
  NAND2X1 gate2675 ( .A(N9368), .B(N9367), .Y(N9702) );
  OR2X1 gate2676 ( .A(N8996), .B(N8517), .Y(N9707) );
  INVX1 gate2677 ( .A(N9183), .Y(N9710) );
  INVX1 gate2678 ( .A(N8996), .Y(N9711) );
  INVX1 gate2679 ( .A(N9193), .Y(N9714) );
  INVX1 gate2680 ( .A(N9203), .Y(N9715) );
  NAND2X1 gate2681 ( .A(N9203), .B(N6235), .Y(N9716) );
  OR2X1 gate2682 ( .A(N9005), .B(N8518), .Y(N9717) );
  INVX1 gate2683 ( .A(N9206), .Y(N9720) );
  INVX1 gate2684 ( .A(N9220), .Y(N9721) );
  NAND2X1 gate2685 ( .A(N9220), .B(N7573), .Y(N9722) );
  INVX1 gate2686 ( .A(N9005), .Y(N9723) );
  INVX1 gate2687 ( .A(N9223), .Y(N9726) );
  NAND2X1 gate2688 ( .A(N9418), .B(N9417), .Y(N9727) );
  AND2X1 gate2689 ( .A(N9268), .B(N8269), .Y(N9732) );
  NAND2X1 gate2690 ( .A(N9581), .B(N9326), .Y(N9733) );
  AND2X1 gate2691_1 ( .A(N89), .B(N9408), .Y(N9734_1) );
  AND2X1 gate2691_2 ( .A(N9332), .B(N8394), .Y(N9734_2) );
  AND2X1 gate2691_3 ( .A(N8421), .B(N9734_1), .Y(N9734_3) );
  AND2X1 gate2691 ( .A(N9734_2), .B(N9734_3), .Y(N9734) );
  AND2X1 gate2692_1 ( .A(N89), .B(N9408), .Y(N9735_1) );
  AND2X1 gate2692_2 ( .A(N9332), .B(N8394), .Y(N9735_2) );
  AND2X1 gate2692_3 ( .A(N8421), .B(N9735_1), .Y(N9735_3) );
  AND2X1 gate2692 ( .A(N9735_2), .B(N9735_3), .Y(N9735) );
  AND2X1 gate2693 ( .A(N9265), .B(N8262), .Y(N9736) );
  INVX1 gate2694 ( .A(N9555), .Y(N9737) );
  INVX1 gate2695 ( .A(N9556), .Y(N9738) );
  NAND2X1 gate2696 ( .A(N9361), .B(N9601), .Y(N9739) );
  NAND2X1 gate2697 ( .A(N9423), .B(N1115), .Y(N9740) );
  INVX1 gate2698 ( .A(N9423), .Y(N9741) );
  NAND2X1 gate2699 ( .A(N9299), .B(N9570), .Y(N9742) );
  AND2X1 gate2700 ( .A(N8333), .B(N9280), .Y(N9754) );
  OR2X1 gate2701 ( .A(N8898), .B(N9560), .Y(N9758) );
  NAND2X1 gate2702 ( .A(N8660), .B(N9561), .Y(N9762) );
  NAND2X1 gate2703 ( .A(N8663), .B(N9563), .Y(N9763) );
  NAND2X1 gate2704 ( .A(N8666), .B(N9565), .Y(N9764) );
  NAND2X1 gate2705 ( .A(N8669), .B(N9567), .Y(N9765) );
  NAND2X1 gate2706 ( .A(N9297), .B(N9569), .Y(N9766) );
  AND2X1 gate2707 ( .A(N9280), .B(N367), .Y(N9767) );
  NAND2X1 gate2708 ( .A(N9557), .B(N9276), .Y(N9768) );
  INVX1 gate2709 ( .A(N9307), .Y(N9769) );
  NAND2X1 gate2710 ( .A(N9307), .B(N367), .Y(N9773) );
  NAND2X1 gate2711 ( .A(N9571), .B(N9301), .Y(N9774) );
  AND2X1 gate2712 ( .A(N8365), .B(N9307), .Y(N9775) );
  OR2X1 gate2713 ( .A(N8920), .B(N9579), .Y(N9779) );
  INVX1 gate2714 ( .A(N9478), .Y(N9784) );
  NAND2X1 gate2715 ( .A(N9616), .B(N9402), .Y(N9785) );
  OR2X1 gate2716 ( .A(N8950), .B(N9585), .Y(N9786) );
  AND2X1 gate2717_1 ( .A(N89), .B(N9408), .Y(N9790_1) );
  AND2X1 gate2717_2 ( .A(N9332), .B(N8394), .Y(N9790_2) );
  AND2X1 gate2717 ( .A(N9790_1), .B(N9790_2), .Y(N9790) );
  OR2X1 gate2718 ( .A(N8963), .B(N9591), .Y(N9791) );
  NAND2X1 gate2719 ( .A(N8735), .B(N9592), .Y(N9795) );
  NAND2X1 gate2720 ( .A(N8738), .B(N9594), .Y(N9796) );
  NAND2X1 gate2721 ( .A(N8741), .B(N9596), .Y(N9797) );
  NAND2X1 gate2722 ( .A(N8744), .B(N9598), .Y(N9798) );
  NAND2X1 gate2723 ( .A(N9359), .B(N9600), .Y(N9799) );
  NOR2X1 gate2724 ( .A(N9602), .B(N9369), .Y(N9800) );
  NOR2X1 gate2725 ( .A(N9603), .B(N9370), .Y(N9801) );
  NOR2X1 gate2726 ( .A(N9604), .B(N9371), .Y(N9802) );
  NOR2X1 gate2727 ( .A(N9605), .B(N9372), .Y(N9803) );
  INVX1 gate2728 ( .A(N9485), .Y(N9805) );
  INVX1 gate2729 ( .A(N9488), .Y(N9806) );
  OR2X1 gate2730 ( .A(N8995), .B(N9611), .Y(N9809) );
  NOR2X1 gate2731 ( .A(N9612), .B(N9396), .Y(N9813) );
  NOR2X1 gate2732 ( .A(N9613), .B(N9397), .Y(N9814) );
  NOR2X1 gate2733 ( .A(N9614), .B(N9398), .Y(N9815) );
  NOR2X1 gate2734 ( .A(N9615), .B(N9399), .Y(N9816) );
  AND2X1 gate2735 ( .A(N9617), .B(N9407), .Y(N9817) );
  OR2X1 gate2736 ( .A(N9029), .B(N9618), .Y(N9820) );
  INVX1 gate2737 ( .A(N9517), .Y(N9825) );
  INVX1 gate2738 ( .A(N9520), .Y(N9826) );
  NOR2X1 gate2739 ( .A(N9621), .B(N9419), .Y(N9827) );
  NOR2X1 gate2740 ( .A(N9622), .B(N9420), .Y(N9828) );
  NOR2X1 gate2741 ( .A(N9623), .B(N9421), .Y(N9829) );
  NOR2X1 gate2742 ( .A(N9624), .B(N9422), .Y(N9830) );
  INVX1 gate2743 ( .A(N9426), .Y(N9835) );
  NAND2X1 gate2744 ( .A(N9426), .B(N4789), .Y(N9836) );
  INVX1 gate2745 ( .A(N9429), .Y(N9837) );
  NAND2X1 gate2746 ( .A(N9429), .B(N4794), .Y(N9838) );
  NAND2X1 gate2747 ( .A(N3625), .B(N9659), .Y(N9846) );
  NAND2X1 gate2748 ( .A(N4810), .B(N9661), .Y(N9847) );
  INVX1 gate2749 ( .A(N9462), .Y(N9862) );
  NAND2X1 gate2750 ( .A(N7553), .B(N9690), .Y(N9863) );
  INVX1 gate2751 ( .A(N9473), .Y(N9866) );
  NAND2X1 gate2752 ( .A(N5030), .B(N9715), .Y(N9873) );
  NAND2X1 gate2753 ( .A(N6236), .B(N9721), .Y(N9876) );
  NAND2X1 gate2754 ( .A(N9795), .B(N9593), .Y(N9890) );
  NAND2X1 gate2755 ( .A(N9797), .B(N9597), .Y(N9891) );
  INVX1 gate2756 ( .A(N9799), .Y(N9892) );
  NAND2X1 gate2757 ( .A(N871), .B(N9741), .Y(N9893) );
  NAND2X1 gate2758 ( .A(N9762), .B(N9562), .Y(N9894) );
  NAND2X1 gate2759 ( .A(N9764), .B(N9566), .Y(N9895) );
  INVX1 gate2760 ( .A(N9766), .Y(N9896) );
  INVX1 gate2761 ( .A(N9626), .Y(N9897) );
  NAND2X1 gate2762 ( .A(N9626), .B(N9249), .Y(N9898) );
  INVX1 gate2763 ( .A(N9629), .Y(N9899) );
  NAND2X1 gate2764 ( .A(N9629), .B(N9250), .Y(N9900) );
  INVX1 gate2765 ( .A(N9632), .Y(N9901) );
  NAND2X1 gate2766 ( .A(N9632), .B(N9251), .Y(N9902) );
  INVX1 gate2767 ( .A(N9635), .Y(N9903) );
  NAND2X1 gate2768 ( .A(N9635), .B(N9252), .Y(N9904) );
  INVX1 gate2769 ( .A(N9543), .Y(N9905) );
  INVX1 gate2770 ( .A(N9650), .Y(N9906) );
  NAND2X1 gate2771 ( .A(N9650), .B(N5769), .Y(N9907) );
  INVX1 gate2772 ( .A(N9653), .Y(N9908) );
  NAND2X1 gate2773 ( .A(N9653), .B(N5770), .Y(N9909) );
  INVX1 gate2774 ( .A(N9656), .Y(N9910) );
  NAND2X1 gate2775 ( .A(N9656), .B(N9262), .Y(N9911) );
  INVX1 gate2776 ( .A(N9551), .Y(N9917) );
  NAND2X1 gate2777 ( .A(N9763), .B(N9564), .Y(N9923) );
  NAND2X1 gate2778 ( .A(N9765), .B(N9568), .Y(N9924) );
  OR2X1 gate2779 ( .A(N8902), .B(N9767), .Y(N9925) );
  AND2X1 gate2780 ( .A(N9575), .B(N9773), .Y(N9932) );
  AND2X1 gate2781 ( .A(N9575), .B(N9769), .Y(N9935) );
  INVX1 gate2782 ( .A(N9698), .Y(N9938) );
  NAND2X1 gate2783 ( .A(N9698), .B(N9323), .Y(N9939) );
  NAND2X1 gate2784 ( .A(N9796), .B(N9595), .Y(N9945) );
  NAND2X1 gate2785 ( .A(N9798), .B(N9599), .Y(N9946) );
  INVX1 gate2786 ( .A(N9702), .Y(N9947) );
  NAND2X1 gate2787 ( .A(N9702), .B(N6102), .Y(N9948) );
  AND2X1 gate2788 ( .A(N9608), .B(N9375), .Y(N9949) );
  INVX1 gate2789 ( .A(N9727), .Y(N9953) );
  NAND2X1 gate2790 ( .A(N9727), .B(N9412), .Y(N9954) );
  NAND2X1 gate2791 ( .A(N3502), .B(N9835), .Y(N9955) );
  NAND2X1 gate2792 ( .A(N3510), .B(N9837), .Y(N9956) );
  INVX1 gate2793 ( .A(N9642), .Y(N9957) );
  NAND2X1 gate2794 ( .A(N9642), .B(N9645), .Y(N9958) );
  INVX1 gate2795 ( .A(N9646), .Y(N9959) );
  NAND2X1 gate2796 ( .A(N9646), .B(N9649), .Y(N9960) );
  NAND2X1 gate2797 ( .A(N9660), .B(N9846), .Y(N9961) );
  NAND2X1 gate2798 ( .A(N9662), .B(N9847), .Y(N9964) );
  INVX1 gate2799 ( .A(N9663), .Y(N9967) );
  NAND2X1 gate2800 ( .A(N9663), .B(N9666), .Y(N9968) );
  INVX1 gate2801 ( .A(N9667), .Y(N9969) );
  NAND2X1 gate2802 ( .A(N9667), .B(N9670), .Y(N9970) );
  INVX1 gate2803 ( .A(N9671), .Y(N9971) );
  NAND2X1 gate2804 ( .A(N9671), .B(N6213), .Y(N9972) );
  INVX1 gate2805 ( .A(N9675), .Y(N9973) );
  NAND2X1 gate2806 ( .A(N9675), .B(N7551), .Y(N9974) );
  INVX1 gate2807 ( .A(N9679), .Y(N9975) );
  NAND2X1 gate2808 ( .A(N9679), .B(N7552), .Y(N9976) );
  INVX1 gate2809 ( .A(N9682), .Y(N9977) );
  INVX1 gate2810 ( .A(N9685), .Y(N9978) );
  NAND2X1 gate2811 ( .A(N9691), .B(N9863), .Y(N9979) );
  INVX1 gate2812 ( .A(N9692), .Y(N9982) );
  NAND2X1 gate2813 ( .A(N9814), .B(N9813), .Y(N9983) );
  NAND2X1 gate2814 ( .A(N9816), .B(N9815), .Y(N9986) );
  NAND2X1 gate2815 ( .A(N9801), .B(N9800), .Y(N9989) );
  NAND2X1 gate2816 ( .A(N9803), .B(N9802), .Y(N9992) );
  INVX1 gate2817 ( .A(N9707), .Y(N9995) );
  NAND2X1 gate2818 ( .A(N9707), .B(N6231), .Y(N9996) );
  INVX1 gate2819 ( .A(N9711), .Y(N9997) );
  NAND2X1 gate2820 ( .A(N9711), .B(N7572), .Y(N9998) );
  NAND2X1 gate2821 ( .A(N9716), .B(N9873), .Y(N9999) );
  INVX1 gate2822 ( .A(N9717), .Y(N10002) );
  NAND2X1 gate2823 ( .A(N9722), .B(N9876), .Y(N10003) );
  INVX1 gate2824 ( .A(N9723), .Y(N10006) );
  NAND2X1 gate2825 ( .A(N9830), .B(N9829), .Y(N10007) );
  NAND2X1 gate2826 ( .A(N9828), .B(N9827), .Y(N10010) );
  AND2X1 gate2827_1 ( .A(N9791), .B(N8307), .Y(N10013_1) );
  AND2X1 gate2827 ( .A(N8269), .B(N10013_1), .Y(N10013) );
  AND2X1 gate2828_1 ( .A(N9758), .B(N9344), .Y(N10014_1) );
  AND2X1 gate2828_2 ( .A(N8307), .B(N8269), .Y(N10014_2) );
  AND2X1 gate2828 ( .A(N10014_1), .B(N10014_2), .Y(N10014) );
  AND2X1 gate2829_1 ( .A(N367), .B(N9754), .Y(N10015_1) );
  AND2X1 gate2829_2 ( .A(N9344), .B(N8307), .Y(N10015_2) );
  AND2X1 gate2829_3 ( .A(N8269), .B(N10015_1), .Y(N10015_3) );
  AND2X1 gate2829 ( .A(N10015_2), .B(N10015_3), .Y(N10015) );
  AND2X1 gate2830_1 ( .A(N9786), .B(N8394), .Y(N10016_1) );
  AND2X1 gate2830 ( .A(N8421), .B(N10016_1), .Y(N10016) );
  AND2X1 gate2831_1 ( .A(N9820), .B(N9332), .Y(N10017_1) );
  AND2X1 gate2831_2 ( .A(N8394), .B(N8421), .Y(N10017_2) );
  AND2X1 gate2831 ( .A(N10017_1), .B(N10017_2), .Y(N10017) );
  AND2X1 gate2832_1 ( .A(N9786), .B(N8394), .Y(N10018_1) );
  AND2X1 gate2832 ( .A(N8421), .B(N10018_1), .Y(N10018) );
  AND2X1 gate2833_1 ( .A(N9820), .B(N9332), .Y(N10019_1) );
  AND2X1 gate2833_2 ( .A(N8394), .B(N8421), .Y(N10019_2) );
  AND2X1 gate2833 ( .A(N10019_1), .B(N10019_2), .Y(N10019) );
  AND2X1 gate2834_1 ( .A(N9809), .B(N8298), .Y(N10020_1) );
  AND2X1 gate2834 ( .A(N8262), .B(N10020_1), .Y(N10020) );
  AND2X1 gate2835_1 ( .A(N9779), .B(N9385), .Y(N10021_1) );
  AND2X1 gate2835_2 ( .A(N8298), .B(N8262), .Y(N10021_2) );
  AND2X1 gate2835 ( .A(N10021_1), .B(N10021_2), .Y(N10021) );
  AND2X1 gate2836_1 ( .A(N367), .B(N9775), .Y(N10022_1) );
  AND2X1 gate2836_2 ( .A(N9385), .B(N8298), .Y(N10022_2) );
  AND2X1 gate2836_3 ( .A(N8262), .B(N10022_1), .Y(N10022_3) );
  AND2X1 gate2836 ( .A(N10022_2), .B(N10022_3), .Y(N10022) );
  INVX1 gate2837 ( .A(N9945), .Y(N10023) );
  INVX1 gate2838 ( .A(N9946), .Y(N10024) );
  NAND2X1 gate2839 ( .A(N9740), .B(N9893), .Y(N10025) );
  INVX1 gate2840 ( .A(N9923), .Y(N10026) );
  INVX1 gate2841 ( .A(N9924), .Y(N10028) );
  NAND2X1 gate2842 ( .A(N8595), .B(N9897), .Y(N10032) );
  NAND2X1 gate2843 ( .A(N8598), .B(N9899), .Y(N10033) );
  NAND2X1 gate2844 ( .A(N8601), .B(N9901), .Y(N10034) );
  NAND2X1 gate2845 ( .A(N8604), .B(N9903), .Y(N10035) );
  NAND2X1 gate2846 ( .A(N4803), .B(N9906), .Y(N10036) );
  NAND2X1 gate2847 ( .A(N4806), .B(N9908), .Y(N10037) );
  NAND2X1 gate2848 ( .A(N8627), .B(N9910), .Y(N10038) );
  AND2X1 gate2849 ( .A(N9809), .B(N8298), .Y(N10039) );
  AND2X1 gate2850_1 ( .A(N9779), .B(N9385), .Y(N10040_1) );
  AND2X1 gate2850 ( .A(N8298), .B(N10040_1), .Y(N10040) );
  AND2X1 gate2851_1 ( .A(N367), .B(N9775), .Y(N10041_1) );
  AND2X1 gate2851_2 ( .A(N9385), .B(N8298), .Y(N10041_2) );
  AND2X1 gate2851 ( .A(N10041_1), .B(N10041_2), .Y(N10041) );
  AND2X1 gate2852 ( .A(N9779), .B(N9385), .Y(N10042) );
  AND2X1 gate2853_1 ( .A(N367), .B(N9775), .Y(N10043_1) );
  AND2X1 gate2853 ( .A(N9385), .B(N10043_1), .Y(N10043) );
  NAND2X1 gate2854 ( .A(N8727), .B(N9938), .Y(N10050) );
  INVX1 gate2855 ( .A(N9817), .Y(N10053) );
  AND2X1 gate2856 ( .A(N9817), .B(N9029), .Y(N10054) );
  AND2X1 gate2857 ( .A(N9786), .B(N8394), .Y(N10055) );
  AND2X1 gate2858_1 ( .A(N9820), .B(N9332), .Y(N10056_1) );
  AND2X1 gate2858 ( .A(N8394), .B(N10056_1), .Y(N10056) );
  AND2X1 gate2859 ( .A(N9791), .B(N8307), .Y(N10057) );
  AND2X1 gate2860_1 ( .A(N9758), .B(N9344), .Y(N10058_1) );
  AND2X1 gate2860 ( .A(N8307), .B(N10058_1), .Y(N10058) );
  AND2X1 gate2861_1 ( .A(N367), .B(N9754), .Y(N10059_1) );
  AND2X1 gate2861_2 ( .A(N9344), .B(N8307), .Y(N10059_2) );
  AND2X1 gate2861 ( .A(N10059_1), .B(N10059_2), .Y(N10059) );
  AND2X1 gate2862 ( .A(N9758), .B(N9344), .Y(N10060) );
  AND2X1 gate2863_1 ( .A(N367), .B(N9754), .Y(N10061_1) );
  AND2X1 gate2863 ( .A(N9344), .B(N10061_1), .Y(N10061) );
  NAND2X1 gate2864 ( .A(N4997), .B(N9947), .Y(N10062) );
  NAND2X1 gate2865 ( .A(N8811), .B(N9953), .Y(N10067) );
  NAND2X1 gate2866 ( .A(N9955), .B(N9836), .Y(N10070) );
  NAND2X1 gate2867 ( .A(N9956), .B(N9838), .Y(N10073) );
  NAND2X1 gate2868 ( .A(N9068), .B(N9957), .Y(N10076) );
  NAND2X1 gate2869 ( .A(N9074), .B(N9959), .Y(N10077) );
  NAND2X1 gate2870 ( .A(N9089), .B(N9967), .Y(N10082) );
  NAND2X1 gate2871 ( .A(N9095), .B(N9969), .Y(N10083) );
  NAND2X1 gate2872 ( .A(N4871), .B(N9971), .Y(N10084) );
  NAND2X1 gate2873 ( .A(N6214), .B(N9973), .Y(N10085) );
  NAND2X1 gate2874 ( .A(N6217), .B(N9975), .Y(N10086) );
  NAND2X1 gate2875 ( .A(N5027), .B(N9995), .Y(N10093) );
  NAND2X1 gate2876 ( .A(N6232), .B(N9997), .Y(N10094) );
  OR2X1 gate2877_1 ( .A(N9238), .B(N9732), .Y(N10101_1) );
  OR2X1 gate2877_2 ( .A(N10013), .B(N10014), .Y(N10101_2) );
  OR2X1 gate2877_3 ( .A(N10015), .B(N10101_1), .Y(N10101_3) );
  OR2X1 gate2877 ( .A(N10101_2), .B(N10101_3), .Y(N10101) );
  OR2X1 gate2878_1 ( .A(N9339), .B(N9526), .Y(N10102_1) );
  OR2X1 gate2878_2 ( .A(N10016), .B(N10017), .Y(N10102_2) );
  OR2X1 gate2878_3 ( .A(N9734), .B(N10102_1), .Y(N10102_3) );
  OR2X1 gate2878 ( .A(N10102_2), .B(N10102_3), .Y(N10102) );
  OR2X1 gate2879_1 ( .A(N9339), .B(N9531), .Y(N10103_1) );
  OR2X1 gate2879_2 ( .A(N10018), .B(N10019), .Y(N10103_2) );
  OR2X1 gate2879_3 ( .A(N9735), .B(N10103_1), .Y(N10103_3) );
  OR2X1 gate2879 ( .A(N10103_2), .B(N10103_3), .Y(N10103) );
  OR2X1 gate2880_1 ( .A(N9242), .B(N9736), .Y(N10104_1) );
  OR2X1 gate2880_2 ( .A(N10020), .B(N10021), .Y(N10104_2) );
  OR2X1 gate2880_3 ( .A(N10022), .B(N10104_1), .Y(N10104_3) );
  OR2X1 gate2880 ( .A(N10104_2), .B(N10104_3), .Y(N10104) );
  AND2X1 gate2881 ( .A(N9925), .B(N9894), .Y(N10105) );
  AND2X1 gate2882 ( .A(N9925), .B(N9895), .Y(N10106) );
  AND2X1 gate2883 ( .A(N9925), .B(N9896), .Y(N10107) );
  AND2X1 gate2884 ( .A(N9925), .B(N8253), .Y(N10108) );
  NAND2X1 gate2885 ( .A(N10032), .B(N9898), .Y(N10109) );
  NAND2X1 gate2886 ( .A(N10033), .B(N9900), .Y(N10110) );
  NAND2X1 gate2887 ( .A(N10034), .B(N9902), .Y(N10111) );
  NAND2X1 gate2888 ( .A(N10035), .B(N9904), .Y(N10112) );
  NAND2X1 gate2889 ( .A(N10036), .B(N9907), .Y(N10113) );
  NAND2X1 gate2890 ( .A(N10037), .B(N9909), .Y(N10114) );
  NAND2X1 gate2891 ( .A(N10038), .B(N9911), .Y(N10115) );
  OR2X1 gate2892_1 ( .A(N9265), .B(N10039), .Y(N10116_1) );
  OR2X1 gate2892_2 ( .A(N10040), .B(N10041), .Y(N10116_2) );
  OR2X1 gate2892 ( .A(N10116_1), .B(N10116_2), .Y(N10116) );
  OR2X1 gate2893_1 ( .A(N9809), .B(N10042), .Y(N10119_1) );
  OR2X1 gate2893 ( .A(N10043), .B(N10119_1), .Y(N10119) );
  INVX1 gate2894 ( .A(N9925), .Y(N10124) );
  AND2X1 gate2895 ( .A(N9768), .B(N9925), .Y(N10130) );
  INVX1 gate2896 ( .A(N9932), .Y(N10131) );
  INVX1 gate2897 ( .A(N9935), .Y(N10132) );
  AND2X1 gate2898 ( .A(N9932), .B(N8920), .Y(N10133) );
  NAND2X1 gate2899 ( .A(N10050), .B(N9939), .Y(N10134) );
  INVX1 gate2900 ( .A(N9983), .Y(N10135) );
  NAND2X1 gate2901 ( .A(N9983), .B(N9324), .Y(N10136) );
  INVX1 gate2902 ( .A(N9986), .Y(N10137) );
  NAND2X1 gate2903 ( .A(N9986), .B(N9784), .Y(N10138) );
  AND2X1 gate2904 ( .A(N9785), .B(N10053), .Y(N10139) );
  OR2X1 gate2905_1 ( .A(N8943), .B(N10055), .Y(N10140_1) );
  OR2X1 gate2905_2 ( .A(N10056), .B(N9790), .Y(N10140_2) );
  OR2X1 gate2905 ( .A(N10140_1), .B(N10140_2), .Y(N10140) );
  OR2X1 gate2906_1 ( .A(N9268), .B(N10057), .Y(N10141_1) );
  OR2X1 gate2906_2 ( .A(N10058), .B(N10059), .Y(N10141_2) );
  OR2X1 gate2906 ( .A(N10141_1), .B(N10141_2), .Y(N10141) );
  OR2X1 gate2907_1 ( .A(N9791), .B(N10060), .Y(N10148_1) );
  OR2X1 gate2907 ( .A(N10061), .B(N10148_1), .Y(N10148) );
  NAND2X1 gate2908 ( .A(N10062), .B(N9948), .Y(N10155) );
  INVX1 gate2909 ( .A(N9989), .Y(N10156) );
  NAND2X1 gate2910 ( .A(N9989), .B(N9805), .Y(N10157) );
  INVX1 gate2911 ( .A(N9992), .Y(N10158) );
  NAND2X1 gate2912 ( .A(N9992), .B(N9806), .Y(N10159) );
  INVX1 gate2913 ( .A(N9949), .Y(N10160) );
  NAND2X1 gate2914 ( .A(N10067), .B(N9954), .Y(N10161) );
  INVX1 gate2915 ( .A(N10007), .Y(N10162) );
  NAND2X1 gate2916 ( .A(N10007), .B(N9825), .Y(N10163) );
  INVX1 gate2917 ( .A(N10010), .Y(N10164) );
  NAND2X1 gate2918 ( .A(N10010), .B(N9826), .Y(N10165) );
  NAND2X1 gate2919 ( .A(N10076), .B(N9958), .Y(N10170) );
  NAND2X1 gate2920 ( .A(N10077), .B(N9960), .Y(N10173) );
  INVX1 gate2921 ( .A(N9961), .Y(N10176) );
  NAND2X1 gate2922 ( .A(N9961), .B(N9082), .Y(N10177) );
  INVX1 gate2923 ( .A(N9964), .Y(N10178) );
  NAND2X1 gate2924 ( .A(N9964), .B(N9086), .Y(N10179) );
  NAND2X1 gate2925 ( .A(N10082), .B(N9968), .Y(N10180) );
  NAND2X1 gate2926 ( .A(N10083), .B(N9970), .Y(N10183) );
  NAND2X1 gate2927 ( .A(N9972), .B(N10084), .Y(N10186) );
  NAND2X1 gate2928 ( .A(N9974), .B(N10085), .Y(N10189) );
  NAND2X1 gate2929 ( .A(N9976), .B(N10086), .Y(N10192) );
  INVX1 gate2930 ( .A(N9979), .Y(N10195) );
  NAND2X1 gate2931 ( .A(N9979), .B(N9982), .Y(N10196) );
  NAND2X1 gate2932 ( .A(N9996), .B(N10093), .Y(N10197) );
  NAND2X1 gate2933 ( .A(N9998), .B(N10094), .Y(N10200) );
  INVX1 gate2934 ( .A(N9999), .Y(N10203) );
  NAND2X1 gate2935 ( .A(N9999), .B(N10002), .Y(N10204) );
  INVX1 gate2936 ( .A(N10003), .Y(N10205) );
  NAND2X1 gate2937 ( .A(N10003), .B(N10006), .Y(N10206) );
  NAND2X1 gate2938 ( .A(N10070), .B(N4308), .Y(N10212) );
  NAND2X1 gate2939 ( .A(N10073), .B(N4313), .Y(N10213) );
  AND2X1 gate2940 ( .A(N9774), .B(N10131), .Y(N10230) );
  NAND2X1 gate2941 ( .A(N8730), .B(N10135), .Y(N10231) );
  NAND2X1 gate2942 ( .A(N9478), .B(N10137), .Y(N10232) );
  OR2X1 gate2943 ( .A(N10139), .B(N10054), .Y(N10233) );
  NAND2X1 gate2944 ( .A(N7100), .B(N10140), .Y(N10234) );
  NAND2X1 gate2945 ( .A(N9485), .B(N10156), .Y(N10237) );
  NAND2X1 gate2946 ( .A(N9488), .B(N10158), .Y(N10238) );
  NAND2X1 gate2947 ( .A(N9517), .B(N10162), .Y(N10239) );
  NAND2X1 gate2948 ( .A(N9520), .B(N10164), .Y(N10240) );
  INVX1 gate2949 ( .A(N10070), .Y(N10241) );
  INVX1 gate2950 ( .A(N10073), .Y(N10242) );
  NAND2X1 gate2951 ( .A(N8146), .B(N10176), .Y(N10247) );
  NAND2X1 gate2952 ( .A(N8156), .B(N10178), .Y(N10248) );
  NAND2X1 gate2953 ( .A(N9692), .B(N10195), .Y(N10259) );
  NAND2X1 gate2954 ( .A(N9717), .B(N10203), .Y(N10264) );
  NAND2X1 gate2955 ( .A(N9723), .B(N10205), .Y(N10265) );
  AND2X1 gate2956 ( .A(N10026), .B(N10124), .Y(N10266) );
  AND2X1 gate2957 ( .A(N10028), .B(N10124), .Y(N10267) );
  AND2X1 gate2958 ( .A(N9742), .B(N10124), .Y(N10268) );
  AND2X1 gate2959 ( .A(N6923), .B(N10124), .Y(N10269) );
  NAND2X1 gate2960 ( .A(N6762), .B(N10116), .Y(N10270) );
  NAND2X1 gate2961 ( .A(N3061), .B(N10241), .Y(N10271) );
  NAND2X1 gate2962 ( .A(N3064), .B(N10242), .Y(N10272) );
  BUFX2 gate2963 ( .A(N10116), .Y(N10273) );
  AND2X1 gate2964_1 ( .A(N10141), .B(N5728), .Y(N10278_1) );
  AND2X1 gate2964_2 ( .A(N5707), .B(N5718), .Y(N10278_2) );
  AND2X1 gate2964_3 ( .A(N5697), .B(N10278_1), .Y(N10278_3) );
  AND2X1 gate2964 ( .A(N10278_2), .B(N10278_3), .Y(N10278) );
  AND2X1 gate2965_1 ( .A(N10141), .B(N5728), .Y(N10279_1) );
  AND2X1 gate2965_2 ( .A(N5707), .B(N5718), .Y(N10279_2) );
  AND2X1 gate2965 ( .A(N10279_1), .B(N10279_2), .Y(N10279) );
  AND2X1 gate2966_1 ( .A(N10141), .B(N5728), .Y(N10280_1) );
  AND2X1 gate2966 ( .A(N5718), .B(N10280_1), .Y(N10280) );
  AND2X1 gate2967 ( .A(N10141), .B(N5728), .Y(N10281) );
  AND2X1 gate2968 ( .A(N6784), .B(N10141), .Y(N10282) );
  INVX1 gate2969 ( .A(N10119), .Y(N10283) );
  AND2X1 gate2970_1 ( .A(N10148), .B(N5936), .Y(N10287_1) );
  AND2X1 gate2970_2 ( .A(N5915), .B(N5926), .Y(N10287_2) );
  AND2X1 gate2970_3 ( .A(N5905), .B(N10287_1), .Y(N10287_3) );
  AND2X1 gate2970 ( .A(N10287_2), .B(N10287_3), .Y(N10287) );
  AND2X1 gate2971_1 ( .A(N10148), .B(N5936), .Y(N10288_1) );
  AND2X1 gate2971_2 ( .A(N5915), .B(N5926), .Y(N10288_2) );
  AND2X1 gate2971 ( .A(N10288_1), .B(N10288_2), .Y(N10288) );
  AND2X1 gate2972_1 ( .A(N10148), .B(N5936), .Y(N10289_1) );
  AND2X1 gate2972 ( .A(N5926), .B(N10289_1), .Y(N10289) );
  AND2X1 gate2973 ( .A(N10148), .B(N5936), .Y(N10290) );
  AND2X1 gate2974 ( .A(N6881), .B(N10148), .Y(N10291) );
  AND2X1 gate2975 ( .A(N8898), .B(N10124), .Y(N10292) );
  NAND2X1 gate2976 ( .A(N10231), .B(N10136), .Y(N10293) );
  NAND2X1 gate2977 ( .A(N10232), .B(N10138), .Y(N10294) );
  NAND2X1 gate2978 ( .A(N8412), .B(N10233), .Y(N10295) );
  AND2X1 gate2979 ( .A(N8959), .B(N10234), .Y(N10296) );
  NAND2X1 gate2980 ( .A(N10237), .B(N10157), .Y(N10299) );
  NAND2X1 gate2981 ( .A(N10238), .B(N10159), .Y(N10300) );
  OR2X1 gate2982 ( .A(N10230), .B(N10133), .Y(N10301) );
  NAND2X1 gate2983 ( .A(N10239), .B(N10163), .Y(N10306) );
  NAND2X1 gate2984 ( .A(N10240), .B(N10165), .Y(N10307) );
  BUFX2 gate2985 ( .A(N10148), .Y(N10308) );
  BUFX2 gate2986 ( .A(N10141), .Y(N10311) );
  INVX1 gate2987 ( .A(N10170), .Y(N10314) );
  NAND2X1 gate2988 ( .A(N10170), .B(N9071), .Y(N10315) );
  INVX1 gate2989 ( .A(N10173), .Y(N10316) );
  NAND2X1 gate2990 ( .A(N10173), .B(N9077), .Y(N10317) );
  NAND2X1 gate2991 ( .A(N10247), .B(N10177), .Y(N10318) );
  NAND2X1 gate2992 ( .A(N10248), .B(N10179), .Y(N10321) );
  INVX1 gate2993 ( .A(N10180), .Y(N10324) );
  NAND2X1 gate2994 ( .A(N10180), .B(N9092), .Y(N10325) );
  INVX1 gate2995 ( .A(N10183), .Y(N10326) );
  NAND2X1 gate2996 ( .A(N10183), .B(N9098), .Y(N10327) );
  INVX1 gate2997 ( .A(N10186), .Y(N10328) );
  NAND2X1 gate2998 ( .A(N10186), .B(N9674), .Y(N10329) );
  INVX1 gate2999 ( .A(N10189), .Y(N10330) );
  NAND2X1 gate3000 ( .A(N10189), .B(N9678), .Y(N10331) );
  INVX1 gate3001 ( .A(N10192), .Y(N10332) );
  NAND2X1 gate3002 ( .A(N10192), .B(N9977), .Y(N10333) );
  NAND2X1 gate3003 ( .A(N10259), .B(N10196), .Y(N10334) );
  INVX1 gate3004 ( .A(N10197), .Y(N10337) );
  NAND2X1 gate3005 ( .A(N10197), .B(N9710), .Y(N10338) );
  INVX1 gate3006 ( .A(N10200), .Y(N10339) );
  NAND2X1 gate3007 ( .A(N10200), .B(N9714), .Y(N10340) );
  NAND2X1 gate3008 ( .A(N10264), .B(N10204), .Y(N10341) );
  NAND2X1 gate3009 ( .A(N10265), .B(N10206), .Y(N10344) );
  OR2X1 gate3010 ( .A(N10266), .B(N10105), .Y(N10350) );
  OR2X1 gate3011 ( .A(N10267), .B(N10106), .Y(N10351) );
  OR2X1 gate3012 ( .A(N10268), .B(N10107), .Y(N10352) );
  OR2X1 gate3013 ( .A(N10269), .B(N10108), .Y(N10353) );
  AND2X1 gate3014 ( .A(N8857), .B(N10270), .Y(N10354) );
  NAND2X1 gate3015 ( .A(N10271), .B(N10212), .Y(N10357) );
  NAND2X1 gate3016 ( .A(N10272), .B(N10213), .Y(N10360) );
  OR2X1 gate3017 ( .A(N7620), .B(N10282), .Y(N10367) );
  OR2X1 gate3018 ( .A(N7671), .B(N10291), .Y(N10375) );
  OR2X1 gate3019 ( .A(N10292), .B(N10130), .Y(N10381) );
  AND2X1 gate3020_1 ( .A(N10114), .B(N10134), .Y(N10388_1) );
  AND2X1 gate3020_2 ( .A(N10293), .B(N10294), .Y(N10388_2) );
  AND2X1 gate3020 ( .A(N10388_1), .B(N10388_2), .Y(N10388) );
  AND2X1 gate3021 ( .A(N9582), .B(N10295), .Y(N10391) );
  AND2X1 gate3022_1 ( .A(N10113), .B(N10115), .Y(N10399_1) );
  AND2X1 gate3022_2 ( .A(N10299), .B(N10300), .Y(N10399_2) );
  AND2X1 gate3022 ( .A(N10399_1), .B(N10399_2), .Y(N10399) );
  AND2X1 gate3023_1 ( .A(N10155), .B(N10161), .Y(N10402_1) );
  AND2X1 gate3023_2 ( .A(N10306), .B(N10307), .Y(N10402_2) );
  AND2X1 gate3023 ( .A(N10402_1), .B(N10402_2), .Y(N10402) );
  OR2X1 gate3024_1 ( .A(N3229), .B(N6888), .Y(N10406_1) );
  OR2X1 gate3024_2 ( .A(N6889), .B(N6890), .Y(N10406_2) );
  OR2X1 gate3024_3 ( .A(N10287), .B(N10406_1), .Y(N10406_3) );
  OR2X1 gate3024 ( .A(N10406_2), .B(N10406_3), .Y(N10406) );
  OR2X1 gate3025_1 ( .A(N3232), .B(N6891), .Y(N10409_1) );
  OR2X1 gate3025_2 ( .A(N6892), .B(N10288), .Y(N10409_2) );
  OR2X1 gate3025 ( .A(N10409_1), .B(N10409_2), .Y(N10409) );
  OR2X1 gate3026_1 ( .A(N3236), .B(N6893), .Y(N10412_1) );
  OR2X1 gate3026 ( .A(N10289), .B(N10412_1), .Y(N10412) );
  OR2X1 gate3027 ( .A(N3241), .B(N10290), .Y(N10415) );
  OR2X1 gate3028_1 ( .A(N3137), .B(N6791), .Y(N10419_1) );
  OR2X1 gate3028_2 ( .A(N6792), .B(N6793), .Y(N10419_2) );
  OR2X1 gate3028_3 ( .A(N10278), .B(N10419_1), .Y(N10419_3) );
  OR2X1 gate3028 ( .A(N10419_2), .B(N10419_3), .Y(N10419) );
  OR2X1 gate3029_1 ( .A(N3140), .B(N6794), .Y(N10422_1) );
  OR2X1 gate3029_2 ( .A(N6795), .B(N10279), .Y(N10422_2) );
  OR2X1 gate3029 ( .A(N10422_1), .B(N10422_2), .Y(N10422) );
  OR2X1 gate3030_1 ( .A(N3144), .B(N6796), .Y(N10425_1) );
  OR2X1 gate3030 ( .A(N10280), .B(N10425_1), .Y(N10425) );
  OR2X1 gate3031 ( .A(N3149), .B(N10281), .Y(N10428) );
  NAND2X1 gate3032 ( .A(N8117), .B(N10314), .Y(N10431) );
  NAND2X1 gate3033 ( .A(N8134), .B(N10316), .Y(N10432) );
  NAND2X1 gate3034 ( .A(N8169), .B(N10324), .Y(N10437) );
  NAND2X1 gate3035 ( .A(N8186), .B(N10326), .Y(N10438) );
  NAND2X1 gate3036 ( .A(N9117), .B(N10328), .Y(N10439) );
  NAND2X1 gate3037 ( .A(N9127), .B(N10330), .Y(N10440) );
  NAND2X1 gate3038 ( .A(N9682), .B(N10332), .Y(N10441) );
  NAND2X1 gate3039 ( .A(N9183), .B(N10337), .Y(N10444) );
  NAND2X1 gate3040 ( .A(N9193), .B(N10339), .Y(N10445) );
  INVX1 gate3041 ( .A(N10296), .Y(N10450) );
  AND2X1 gate3042 ( .A(N10296), .B(N4193), .Y(N10451) );
  INVX1 gate3043 ( .A(N10308), .Y(N10455) );
  NAND2X1 gate3044 ( .A(N10308), .B(N8242), .Y(N10456) );
  INVX1 gate3045 ( .A(N10311), .Y(N10465) );
  NAND2X1 gate3046 ( .A(N10311), .B(N8247), .Y(N10466) );
  INVX1 gate3047 ( .A(N10273), .Y(N10479) );
  INVX1 gate3048 ( .A(N10301), .Y(N10497) );
  NAND2X1 gate3049 ( .A(N10431), .B(N10315), .Y(N10509) );
  NAND2X1 gate3050 ( .A(N10432), .B(N10317), .Y(N10512) );
  INVX1 gate3051 ( .A(N10318), .Y(N10515) );
  NAND2X1 gate3052 ( .A(N10318), .B(N8632), .Y(N10516) );
  INVX1 gate3053 ( .A(N10321), .Y(N10517) );
  NAND2X1 gate3054 ( .A(N10321), .B(N8637), .Y(N10518) );
  NAND2X1 gate3055 ( .A(N10437), .B(N10325), .Y(N10519) );
  NAND2X1 gate3056 ( .A(N10438), .B(N10327), .Y(N10522) );
  NAND2X1 gate3057 ( .A(N10439), .B(N10329), .Y(N10525) );
  NAND2X1 gate3058 ( .A(N10440), .B(N10331), .Y(N10528) );
  NAND2X1 gate3059 ( .A(N10441), .B(N10333), .Y(N10531) );
  INVX1 gate3060 ( .A(N10334), .Y(N10534) );
  NAND2X1 gate3061 ( .A(N10334), .B(N9695), .Y(N10535) );
  NAND2X1 gate3062 ( .A(N10444), .B(N10338), .Y(N10536) );
  NAND2X1 gate3063 ( .A(N10445), .B(N10340), .Y(N10539) );
  INVX1 gate3064 ( .A(N10341), .Y(N10542) );
  NAND2X1 gate3065 ( .A(N10341), .B(N9720), .Y(N10543) );
  INVX1 gate3066 ( .A(N10344), .Y(N10544) );
  NAND2X1 gate3067 ( .A(N10344), .B(N9726), .Y(N10545) );
  AND2X1 gate3068 ( .A(N5631), .B(N10450), .Y(N10546) );
  INVX1 gate3069 ( .A(N10391), .Y(N10547) );
  AND2X1 gate3070 ( .A(N10391), .B(N8950), .Y(N10548) );
  AND2X1 gate3071 ( .A(N5165), .B(N10367), .Y(N10549) );
  INVX1 gate3072 ( .A(N10354), .Y(N10550) );
  AND2X1 gate3073 ( .A(N10354), .B(N3126), .Y(N10551) );
  NAND2X1 gate3074 ( .A(N7411), .B(N10455), .Y(N10552) );
  AND2X1 gate3075 ( .A(N10375), .B(N9539), .Y(N10553) );
  AND2X1 gate3076 ( .A(N10375), .B(N9540), .Y(N10554) );
  AND2X1 gate3077 ( .A(N10375), .B(N9541), .Y(N10555) );
  AND2X1 gate3078 ( .A(N10375), .B(N6761), .Y(N10556) );
  INVX1 gate3079 ( .A(N10406), .Y(N10557) );
  NAND2X1 gate3080 ( .A(N10406), .B(N8243), .Y(N10558) );
  INVX1 gate3081 ( .A(N10409), .Y(N10559) );
  NAND2X1 gate3082 ( .A(N10409), .B(N8244), .Y(N10560) );
  INVX1 gate3083 ( .A(N10412), .Y(N10561) );
  NAND2X1 gate3084 ( .A(N10412), .B(N8245), .Y(N10562) );
  INVX1 gate3085 ( .A(N10415), .Y(N10563) );
  NAND2X1 gate3086 ( .A(N10415), .B(N8246), .Y(N10564) );
  NAND2X1 gate3087 ( .A(N7426), .B(N10465), .Y(N10565) );
  INVX1 gate3088 ( .A(N10419), .Y(N10566) );
  NAND2X1 gate3089 ( .A(N10419), .B(N8248), .Y(N10567) );
  INVX1 gate3090 ( .A(N10422), .Y(N10568) );
  NAND2X1 gate3091 ( .A(N10422), .B(N8249), .Y(N10569) );
  INVX1 gate3092 ( .A(N10425), .Y(N10570) );
  NAND2X1 gate3093 ( .A(N10425), .B(N8250), .Y(N10571) );
  INVX1 gate3094 ( .A(N10428), .Y(N10572) );
  NAND2X1 gate3095 ( .A(N10428), .B(N8251), .Y(N10573) );
  INVX1 gate3096 ( .A(N10399), .Y(N10574) );
  INVX1 gate3097 ( .A(N10402), .Y(N10575) );
  INVX1 gate3098 ( .A(N10388), .Y(N10576) );
  AND2X1 gate3099_1 ( .A(N10399), .B(N10402), .Y(N10577_1) );
  AND2X1 gate3099 ( .A(N10388), .B(N10577_1), .Y(N10577) );
  AND2X1 gate3100_1 ( .A(N10360), .B(N9543), .Y(N10581_1) );
  AND2X1 gate3100 ( .A(N10273), .B(N10581_1), .Y(N10581) );
  AND2X1 gate3101_1 ( .A(N10357), .B(N9905), .Y(N10582_1) );
  AND2X1 gate3101 ( .A(N10273), .B(N10582_1), .Y(N10582) );
  INVX1 gate3102 ( .A(N10367), .Y(N10583) );
  AND2X1 gate3103 ( .A(N10367), .B(N5735), .Y(N10587) );
  AND2X1 gate3104 ( .A(N10367), .B(N3135), .Y(N10588) );
  INVX1 gate3105 ( .A(N10375), .Y(N10589) );
  AND2X1 gate3106_1 ( .A(N10381), .B(N7180), .Y(N10594_1) );
  AND2X1 gate3106_2 ( .A(N7159), .B(N7170), .Y(N10594_2) );
  AND2X1 gate3106_3 ( .A(N7149), .B(N10594_1), .Y(N10594_3) );
  AND2X1 gate3106 ( .A(N10594_2), .B(N10594_3), .Y(N10594) );
  AND2X1 gate3107_1 ( .A(N10381), .B(N7180), .Y(N10595_1) );
  AND2X1 gate3107_2 ( .A(N7159), .B(N7170), .Y(N10595_2) );
  AND2X1 gate3107 ( .A(N10595_1), .B(N10595_2), .Y(N10595) );
  AND2X1 gate3108_1 ( .A(N10381), .B(N7180), .Y(N10596_1) );
  AND2X1 gate3108 ( .A(N7170), .B(N10596_1), .Y(N10596) );
  AND2X1 gate3109 ( .A(N10381), .B(N7180), .Y(N10597) );
  AND2X1 gate3110 ( .A(N8444), .B(N10381), .Y(N10598) );
  BUFX2 gate3111 ( .A(N10381), .Y(N10602) );
  NAND2X1 gate3112 ( .A(N7479), .B(N10515), .Y(N10609) );
  NAND2X1 gate3113 ( .A(N7491), .B(N10517), .Y(N10610) );
  NAND2X1 gate3114 ( .A(N9149), .B(N10534), .Y(N10621) );
  NAND2X1 gate3115 ( .A(N9206), .B(N10542), .Y(N10626) );
  NAND2X1 gate3116 ( .A(N9223), .B(N10544), .Y(N10627) );
  OR2X1 gate3117 ( .A(N10546), .B(N10451), .Y(N10628) );
  AND2X1 gate3118 ( .A(N9733), .B(N10547), .Y(N10629) );
  AND2X1 gate3119 ( .A(N5166), .B(N10550), .Y(N10631) );
  NAND2X1 gate3120 ( .A(N10552), .B(N10456), .Y(N10632) );
  NAND2X1 gate3121 ( .A(N7414), .B(N10557), .Y(N10637) );
  NAND2X1 gate3122 ( .A(N7417), .B(N10559), .Y(N10638) );
  NAND2X1 gate3123 ( .A(N7420), .B(N10561), .Y(N10639) );
  NAND2X1 gate3124 ( .A(N7423), .B(N10563), .Y(N10640) );
  NAND2X1 gate3125 ( .A(N10565), .B(N10466), .Y(N10641) );
  NAND2X1 gate3126 ( .A(N7429), .B(N10566), .Y(N10642) );
  NAND2X1 gate3127 ( .A(N7432), .B(N10568), .Y(N10643) );
  NAND2X1 gate3128 ( .A(N7435), .B(N10570), .Y(N10644) );
  NAND2X1 gate3129 ( .A(N7438), .B(N10572), .Y(N10645) );
  AND2X1 gate3130_1 ( .A(N886), .B(N887), .Y(N10647_1) );
  AND2X1 gate3130 ( .A(N10577), .B(N10647_1), .Y(N10647) );
  AND2X1 gate3131_1 ( .A(N10360), .B(N8857), .Y(N10648_1) );
  AND2X1 gate3131 ( .A(N10479), .B(N10648_1), .Y(N10648) );
  AND2X1 gate3132_1 ( .A(N10357), .B(N7609), .Y(N10649_1) );
  AND2X1 gate3132 ( .A(N10479), .B(N10649_1), .Y(N10649) );
  OR2X1 gate3133 ( .A(N8966), .B(N10598), .Y(N10652) );
  OR2X1 gate3134_1 ( .A(N4675), .B(N8451), .Y(N10659_1) );
  OR2X1 gate3134_2 ( .A(N8452), .B(N8453), .Y(N10659_2) );
  OR2X1 gate3134_3 ( .A(N10594), .B(N10659_1), .Y(N10659_3) );
  OR2X1 gate3134 ( .A(N10659_2), .B(N10659_3), .Y(N10659) );
  OR2X1 gate3135_1 ( .A(N4678), .B(N8454), .Y(N10662_1) );
  OR2X1 gate3135_2 ( .A(N8455), .B(N10595), .Y(N10662_2) );
  OR2X1 gate3135 ( .A(N10662_1), .B(N10662_2), .Y(N10662) );
  OR2X1 gate3136_1 ( .A(N4682), .B(N8456), .Y(N10665_1) );
  OR2X1 gate3136 ( .A(N10596), .B(N10665_1), .Y(N10665) );
  OR2X1 gate3137 ( .A(N4687), .B(N10597), .Y(N10668) );
  INVX1 gate3138 ( .A(N10509), .Y(N10671) );
  NAND2X1 gate3139 ( .A(N10509), .B(N8615), .Y(N10672) );
  INVX1 gate3140 ( .A(N10512), .Y(N10673) );
  NAND2X1 gate3141 ( .A(N10512), .B(N8624), .Y(N10674) );
  NAND2X1 gate3142 ( .A(N10609), .B(N10516), .Y(N10675) );
  NAND2X1 gate3143 ( .A(N10610), .B(N10518), .Y(N10678) );
  INVX1 gate3144 ( .A(N10519), .Y(N10681) );
  NAND2X1 gate3145 ( .A(N10519), .B(N8644), .Y(N10682) );
  INVX1 gate3146 ( .A(N10522), .Y(N10683) );
  NAND2X1 gate3147 ( .A(N10522), .B(N8653), .Y(N10684) );
  INVX1 gate3148 ( .A(N10525), .Y(N10685) );
  NAND2X1 gate3149 ( .A(N10525), .B(N9454), .Y(N10686) );
  INVX1 gate3150 ( .A(N10528), .Y(N10687) );
  NAND2X1 gate3151 ( .A(N10528), .B(N9459), .Y(N10688) );
  INVX1 gate3152 ( .A(N10531), .Y(N10689) );
  NAND2X1 gate3153 ( .A(N10531), .B(N9978), .Y(N10690) );
  NAND2X1 gate3154 ( .A(N10621), .B(N10535), .Y(N10691) );
  INVX1 gate3155 ( .A(N10536), .Y(N10694) );
  NAND2X1 gate3156 ( .A(N10536), .B(N9493), .Y(N10695) );
  INVX1 gate3157 ( .A(N10539), .Y(N10696) );
  NAND2X1 gate3158 ( .A(N10539), .B(N9498), .Y(N10697) );
  NAND2X1 gate3159 ( .A(N10626), .B(N10543), .Y(N10698) );
  NAND2X1 gate3160 ( .A(N10627), .B(N10545), .Y(N10701) );
  OR2X1 gate3161 ( .A(N10629), .B(N10548), .Y(N10704) );
  AND2X1 gate3162 ( .A(N3159), .B(N10583), .Y(N10705) );
  OR2X1 gate3163 ( .A(N10631), .B(N10551), .Y(N10706) );
  AND2X1 gate3164 ( .A(N9737), .B(N10589), .Y(N10707) );
  AND2X1 gate3165 ( .A(N9738), .B(N10589), .Y(N10708) );
  AND2X1 gate3166 ( .A(N9243), .B(N10589), .Y(N10709) );
  AND2X1 gate3167 ( .A(N5892), .B(N10589), .Y(N10710) );
  NAND2X1 gate3168 ( .A(N10637), .B(N10558), .Y(N10711) );
  NAND2X1 gate3169 ( .A(N10638), .B(N10560), .Y(N10712) );
  NAND2X1 gate3170 ( .A(N10639), .B(N10562), .Y(N10713) );
  NAND2X1 gate3171 ( .A(N10640), .B(N10564), .Y(N10714) );
  NAND2X1 gate3172 ( .A(N10642), .B(N10567), .Y(N10715) );
  NAND2X1 gate3173 ( .A(N10643), .B(N10569), .Y(N10716) );
  NAND2X1 gate3174 ( .A(N10644), .B(N10571), .Y(N10717) );
  NAND2X1 gate3175 ( .A(N10645), .B(N10573), .Y(N10718) );
  INVX1 gate3176 ( .A(N10602), .Y(N10719) );
  NAND2X1 gate3177 ( .A(N10602), .B(N9244), .Y(N10720) );
  INVX1 gate3178 ( .A(N10647), .Y(N10729) );
  AND2X1 gate3179 ( .A(N5178), .B(N10583), .Y(N10730) );
  AND2X1 gate3180 ( .A(N2533), .B(N10583), .Y(N10731) );
  NAND2X1 gate3181 ( .A(N7447), .B(N10671), .Y(N10737) );
  NAND2X1 gate3182 ( .A(N7465), .B(N10673), .Y(N10738) );
  OR2X1 gate3183_1 ( .A(N10648), .B(N10649), .Y(N10739_1) );
  OR2X1 gate3183_2 ( .A(N10581), .B(N10582), .Y(N10739_2) );
  OR2X1 gate3183 ( .A(N10739_1), .B(N10739_2), .Y(N10739) );
  NAND2X1 gate3184 ( .A(N7503), .B(N10681), .Y(N10746) );
  NAND2X1 gate3185 ( .A(N7521), .B(N10683), .Y(N10747) );
  NAND2X1 gate3186 ( .A(N8678), .B(N10685), .Y(N10748) );
  NAND2X1 gate3187 ( .A(N8690), .B(N10687), .Y(N10749) );
  NAND2X1 gate3188 ( .A(N9685), .B(N10689), .Y(N10750) );
  NAND2X1 gate3189 ( .A(N8757), .B(N10694), .Y(N10753) );
  NAND2X1 gate3190 ( .A(N8769), .B(N10696), .Y(N10754) );
  OR2X1 gate3191 ( .A(N10705), .B(N10549), .Y(N10759) );
  OR2X1 gate3192 ( .A(N10707), .B(N10553), .Y(N10760) );
  OR2X1 gate3193 ( .A(N10708), .B(N10554), .Y(N10761) );
  OR2X1 gate3194 ( .A(N10709), .B(N10555), .Y(N10762) );
  OR2X1 gate3195 ( .A(N10710), .B(N10556), .Y(N10763) );
  NAND2X1 gate3196 ( .A(N8580), .B(N10719), .Y(N10764) );
  AND2X1 gate3197 ( .A(N10652), .B(N9890), .Y(N10765) );
  AND2X1 gate3198 ( .A(N10652), .B(N9891), .Y(N10766) );
  AND2X1 gate3199 ( .A(N10652), .B(N9892), .Y(N10767) );
  AND2X1 gate3200 ( .A(N10652), .B(N8252), .Y(N10768) );
  INVX1 gate3201 ( .A(N10659), .Y(N10769) );
  NAND2X1 gate3202 ( .A(N10659), .B(N9245), .Y(N10770) );
  INVX1 gate3203 ( .A(N10662), .Y(N10771) );
  NAND2X1 gate3204 ( .A(N10662), .B(N9246), .Y(N10772) );
  INVX1 gate3205 ( .A(N10665), .Y(N10773) );
  NAND2X1 gate3206 ( .A(N10665), .B(N9247), .Y(N10774) );
  INVX1 gate3207 ( .A(N10668), .Y(N10775) );
  NAND2X1 gate3208 ( .A(N10668), .B(N9248), .Y(N10776) );
  OR2X1 gate3209 ( .A(N10730), .B(N10587), .Y(N10778) );
  OR2X1 gate3210 ( .A(N10731), .B(N10588), .Y(N10781) );
  INVX1 gate3211 ( .A(N10652), .Y(N10784) );
  NAND2X1 gate3212 ( .A(N10737), .B(N10672), .Y(N10789) );
  NAND2X1 gate3213 ( .A(N10738), .B(N10674), .Y(N10792) );
  INVX1 gate3214 ( .A(N10675), .Y(N10796) );
  NAND2X1 gate3215 ( .A(N10675), .B(N8633), .Y(N10797) );
  INVX1 gate3216 ( .A(N10678), .Y(N10798) );
  NAND2X1 gate3217 ( .A(N10678), .B(N8638), .Y(N10799) );
  NAND2X1 gate3218 ( .A(N10746), .B(N10682), .Y(N10800) );
  NAND2X1 gate3219 ( .A(N10747), .B(N10684), .Y(N10803) );
  NAND2X1 gate3220 ( .A(N10748), .B(N10686), .Y(N10806) );
  NAND2X1 gate3221 ( .A(N10749), .B(N10688), .Y(N10809) );
  NAND2X1 gate3222 ( .A(N10750), .B(N10690), .Y(N10812) );
  INVX1 gate3223 ( .A(N10691), .Y(N10815) );
  NAND2X1 gate3224 ( .A(N10691), .B(N9866), .Y(N10816) );
  NAND2X1 gate3225 ( .A(N10753), .B(N10695), .Y(N10817) );
  NAND2X1 gate3226 ( .A(N10754), .B(N10697), .Y(N10820) );
  INVX1 gate3227 ( .A(N10698), .Y(N10823) );
  NAND2X1 gate3228 ( .A(N10698), .B(N9505), .Y(N10824) );
  INVX1 gate3229 ( .A(N10701), .Y(N10825) );
  NAND2X1 gate3230 ( .A(N10701), .B(N9514), .Y(N10826) );
  NAND2X1 gate3231 ( .A(N10764), .B(N10720), .Y(N10827) );
  NAND2X1 gate3232 ( .A(N8583), .B(N10769), .Y(N10832) );
  NAND2X1 gate3233 ( .A(N8586), .B(N10771), .Y(N10833) );
  NAND2X1 gate3234 ( .A(N8589), .B(N10773), .Y(N10834) );
  NAND2X1 gate3235 ( .A(N8592), .B(N10775), .Y(N10835) );
  INVX1 gate3236 ( .A(N10739), .Y(N10836) );
  BUFX2 gate3237 ( .A(N10778), .Y(N10837) );
  BUFX2 gate3238 ( .A(N10778), .Y(N10838) );
  BUFX2 gate3239 ( .A(N10781), .Y(N10839) );
  BUFX2 gate3240 ( .A(N10781), .Y(N10840) );
  NAND2X1 gate3241 ( .A(N7482), .B(N10796), .Y(N10845) );
  NAND2X1 gate3242 ( .A(N7494), .B(N10798), .Y(N10846) );
  NAND2X1 gate3243 ( .A(N9473), .B(N10815), .Y(N10857) );
  NAND2X1 gate3244 ( .A(N8781), .B(N10823), .Y(N10862) );
  NAND2X1 gate3245 ( .A(N8799), .B(N10825), .Y(N10863) );
  AND2X1 gate3246 ( .A(N10023), .B(N10784), .Y(N10864) );
  AND2X1 gate3247 ( .A(N10024), .B(N10784), .Y(N10865) );
  AND2X1 gate3248 ( .A(N9739), .B(N10784), .Y(N10866) );
  AND2X1 gate3249 ( .A(N7136), .B(N10784), .Y(N10867) );
  NAND2X1 gate3250 ( .A(N10832), .B(N10770), .Y(N10868) );
  NAND2X1 gate3251 ( .A(N10833), .B(N10772), .Y(N10869) );
  NAND2X1 gate3252 ( .A(N10834), .B(N10774), .Y(N10870) );
  NAND2X1 gate3253 ( .A(N10835), .B(N10776), .Y(N10871) );
  INVX1 gate3254 ( .A(N10789), .Y(N10872) );
  NAND2X1 gate3255 ( .A(N10789), .B(N8616), .Y(N10873) );
  INVX1 gate3256 ( .A(N10792), .Y(N10874) );
  NAND2X1 gate3257 ( .A(N10792), .B(N8625), .Y(N10875) );
  NAND2X1 gate3258 ( .A(N10845), .B(N10797), .Y(N10876) );
  NAND2X1 gate3259 ( .A(N10846), .B(N10799), .Y(N10879) );
  INVX1 gate3260 ( .A(N10800), .Y(N10882) );
  NAND2X1 gate3261 ( .A(N10800), .B(N8645), .Y(N10883) );
  INVX1 gate3262 ( .A(N10803), .Y(N10884) );
  NAND2X1 gate3263 ( .A(N10803), .B(N8654), .Y(N10885) );
  INVX1 gate3264 ( .A(N10806), .Y(N10886) );
  NAND2X1 gate3265 ( .A(N10806), .B(N9455), .Y(N10887) );
  INVX1 gate3266 ( .A(N10809), .Y(N10888) );
  NAND2X1 gate3267 ( .A(N10809), .B(N9460), .Y(N10889) );
  INVX1 gate3268 ( .A(N10812), .Y(N10890) );
  NAND2X1 gate3269 ( .A(N10812), .B(N9862), .Y(N10891) );
  NAND2X1 gate3270 ( .A(N10857), .B(N10816), .Y(N10892) );
  INVX1 gate3271 ( .A(N10817), .Y(N10895) );
  NAND2X1 gate3272 ( .A(N10817), .B(N9494), .Y(N10896) );
  INVX1 gate3273 ( .A(N10820), .Y(N10897) );
  NAND2X1 gate3274 ( .A(N10820), .B(N9499), .Y(N10898) );
  NAND2X1 gate3275 ( .A(N10862), .B(N10824), .Y(N10899) );
  NAND2X1 gate3276 ( .A(N10863), .B(N10826), .Y(N10902) );
  OR2X1 gate3277 ( .A(N10864), .B(N10765), .Y(N10905) );
  OR2X1 gate3278 ( .A(N10865), .B(N10766), .Y(N10906) );
  OR2X1 gate3279 ( .A(N10866), .B(N10767), .Y(N10907) );
  OR2X1 gate3280 ( .A(N10867), .B(N10768), .Y(N10908) );
  NAND2X1 gate3281 ( .A(N7450), .B(N10872), .Y(N10909) );
  NAND2X1 gate3282 ( .A(N7468), .B(N10874), .Y(N10910) );
  NAND2X1 gate3283 ( .A(N7506), .B(N10882), .Y(N10915) );
  NAND2X1 gate3284 ( .A(N7524), .B(N10884), .Y(N10916) );
  NAND2X1 gate3285 ( .A(N8681), .B(N10886), .Y(N10917) );
  NAND2X1 gate3286 ( .A(N8693), .B(N10888), .Y(N10918) );
  NAND2X1 gate3287 ( .A(N9462), .B(N10890), .Y(N10919) );
  NAND2X1 gate3288 ( .A(N8760), .B(N10895), .Y(N10922) );
  NAND2X1 gate3289 ( .A(N8772), .B(N10897), .Y(N10923) );
  NAND2X1 gate3290 ( .A(N10909), .B(N10873), .Y(N10928) );
  NAND2X1 gate3291 ( .A(N10910), .B(N10875), .Y(N10931) );
  INVX1 gate3292 ( .A(N10876), .Y(N10934) );
  NAND2X1 gate3293 ( .A(N10876), .B(N8634), .Y(N10935) );
  INVX1 gate3294 ( .A(N10879), .Y(N10936) );
  NAND2X1 gate3295 ( .A(N10879), .B(N8639), .Y(N10937) );
  NAND2X1 gate3296 ( .A(N10915), .B(N10883), .Y(N10938) );
  NAND2X1 gate3297 ( .A(N10916), .B(N10885), .Y(N10941) );
  NAND2X1 gate3298 ( .A(N10917), .B(N10887), .Y(N10944) );
  NAND2X1 gate3299 ( .A(N10918), .B(N10889), .Y(N10947) );
  NAND2X1 gate3300 ( .A(N10919), .B(N10891), .Y(N10950) );
  INVX1 gate3301 ( .A(N10892), .Y(N10953) );
  NAND2X1 gate3302 ( .A(N10892), .B(N9476), .Y(N10954) );
  NAND2X1 gate3303 ( .A(N10922), .B(N10896), .Y(N10955) );
  NAND2X1 gate3304 ( .A(N10923), .B(N10898), .Y(N10958) );
  INVX1 gate3305 ( .A(N10899), .Y(N10961) );
  NAND2X1 gate3306 ( .A(N10899), .B(N9506), .Y(N10962) );
  INVX1 gate3307 ( .A(N10902), .Y(N10963) );
  NAND2X1 gate3308 ( .A(N10902), .B(N9515), .Y(N10964) );
  NAND2X1 gate3309 ( .A(N7485), .B(N10934), .Y(N10969) );
  NAND2X1 gate3310 ( .A(N7497), .B(N10936), .Y(N10970) );
  NAND2X1 gate3311 ( .A(N8718), .B(N10953), .Y(N10981) );
  NAND2X1 gate3312 ( .A(N8784), .B(N10961), .Y(N10986) );
  NAND2X1 gate3313 ( .A(N8802), .B(N10963), .Y(N10987) );
  INVX1 gate3314 ( .A(N10928), .Y(N10988) );
  NAND2X1 gate3315 ( .A(N10928), .B(N8617), .Y(N10989) );
  INVX1 gate3316 ( .A(N10931), .Y(N10990) );
  NAND2X1 gate3317 ( .A(N10931), .B(N8626), .Y(N10991) );
  NAND2X1 gate3318 ( .A(N10969), .B(N10935), .Y(N10992) );
  NAND2X1 gate3319 ( .A(N10970), .B(N10937), .Y(N10995) );
  INVX1 gate3320 ( .A(N10938), .Y(N10998) );
  NAND2X1 gate3321 ( .A(N10938), .B(N8646), .Y(N10999) );
  INVX1 gate3322 ( .A(N10941), .Y(N11000) );
  NAND2X1 gate3323 ( .A(N10941), .B(N8655), .Y(N11001) );
  INVX1 gate3324 ( .A(N10944), .Y(N11002) );
  NAND2X1 gate3325 ( .A(N10944), .B(N9456), .Y(N11003) );
  INVX1 gate3326 ( .A(N10947), .Y(N11004) );
  NAND2X1 gate3327 ( .A(N10947), .B(N9461), .Y(N11005) );
  INVX1 gate3328 ( .A(N10950), .Y(N11006) );
  NAND2X1 gate3329 ( .A(N10950), .B(N9465), .Y(N11007) );
  NAND2X1 gate3330 ( .A(N10981), .B(N10954), .Y(N11008) );
  INVX1 gate3331 ( .A(N10955), .Y(N11011) );
  NAND2X1 gate3332 ( .A(N10955), .B(N9495), .Y(N11012) );
  INVX1 gate3333 ( .A(N10958), .Y(N11013) );
  NAND2X1 gate3334 ( .A(N10958), .B(N9500), .Y(N11014) );
  NAND2X1 gate3335 ( .A(N10986), .B(N10962), .Y(N11015) );
  NAND2X1 gate3336 ( .A(N10987), .B(N10964), .Y(N11018) );
  NAND2X1 gate3337 ( .A(N7453), .B(N10988), .Y(N11023) );
  NAND2X1 gate3338 ( .A(N7471), .B(N10990), .Y(N11024) );
  NAND2X1 gate3339 ( .A(N7509), .B(N10998), .Y(N11027) );
  NAND2X1 gate3340 ( .A(N7527), .B(N11000), .Y(N11028) );
  NAND2X1 gate3341 ( .A(N8684), .B(N11002), .Y(N11029) );
  NAND2X1 gate3342 ( .A(N8696), .B(N11004), .Y(N11030) );
  NAND2X1 gate3343 ( .A(N8702), .B(N11006), .Y(N11031) );
  NAND2X1 gate3344 ( .A(N8763), .B(N11011), .Y(N11034) );
  NAND2X1 gate3345 ( .A(N8775), .B(N11013), .Y(N11035) );
  INVX1 gate3346 ( .A(N10992), .Y(N11040) );
  NAND2X1 gate3347 ( .A(N10992), .B(N8294), .Y(N11041) );
  INVX1 gate3348 ( .A(N10995), .Y(N11042) );
  NAND2X1 gate3349 ( .A(N10995), .B(N8295), .Y(N11043) );
  NAND2X1 gate3350 ( .A(N11023), .B(N10989), .Y(N11044) );
  NAND2X1 gate3351 ( .A(N11024), .B(N10991), .Y(N11047) );
  NAND2X1 gate3352 ( .A(N11027), .B(N10999), .Y(N11050) );
  NAND2X1 gate3353 ( .A(N11028), .B(N11001), .Y(N11053) );
  NAND2X1 gate3354 ( .A(N11029), .B(N11003), .Y(N11056) );
  NAND2X1 gate3355 ( .A(N11030), .B(N11005), .Y(N11059) );
  NAND2X1 gate3356 ( .A(N11031), .B(N11007), .Y(N11062) );
  INVX1 gate3357 ( .A(N11008), .Y(N11065) );
  NAND2X1 gate3358 ( .A(N11008), .B(N9477), .Y(N11066) );
  NAND2X1 gate3359 ( .A(N11034), .B(N11012), .Y(N11067) );
  NAND2X1 gate3360 ( .A(N11035), .B(N11014), .Y(N11070) );
  INVX1 gate3361 ( .A(N11015), .Y(N11073) );
  NAND2X1 gate3362 ( .A(N11015), .B(N9507), .Y(N11074) );
  INVX1 gate3363 ( .A(N11018), .Y(N11075) );
  NAND2X1 gate3364 ( .A(N11018), .B(N9516), .Y(N11076) );
  NAND2X1 gate3365 ( .A(N7488), .B(N11040), .Y(N11077) );
  NAND2X1 gate3366 ( .A(N7500), .B(N11042), .Y(N11078) );
  NAND2X1 gate3367 ( .A(N8721), .B(N11065), .Y(N11095) );
  NAND2X1 gate3368 ( .A(N8787), .B(N11073), .Y(N11098) );
  NAND2X1 gate3369 ( .A(N8805), .B(N11075), .Y(N11099) );
  NAND2X1 gate3370 ( .A(N11077), .B(N11041), .Y(N11100) );
  NAND2X1 gate3371 ( .A(N11078), .B(N11043), .Y(N11103) );
  INVX1 gate3372 ( .A(N11056), .Y(N11106) );
  NAND2X1 gate3373 ( .A(N11056), .B(N9319), .Y(N11107) );
  INVX1 gate3374 ( .A(N11059), .Y(N11108) );
  NAND2X1 gate3375 ( .A(N11059), .B(N9320), .Y(N11109) );
  INVX1 gate3376 ( .A(N11067), .Y(N11110) );
  NAND2X1 gate3377 ( .A(N11067), .B(N9381), .Y(N11111) );
  INVX1 gate3378 ( .A(N11070), .Y(N11112) );
  NAND2X1 gate3379 ( .A(N11070), .B(N9382), .Y(N11113) );
  INVX1 gate3380 ( .A(N11044), .Y(N11114) );
  NAND2X1 gate3381 ( .A(N11044), .B(N8618), .Y(N11115) );
  INVX1 gate3382 ( .A(N11047), .Y(N11116) );
  NAND2X1 gate3383 ( .A(N11047), .B(N8619), .Y(N11117) );
  INVX1 gate3384 ( .A(N11050), .Y(N11118) );
  NAND2X1 gate3385 ( .A(N11050), .B(N8647), .Y(N11119) );
  INVX1 gate3386 ( .A(N11053), .Y(N11120) );
  NAND2X1 gate3387 ( .A(N11053), .B(N8648), .Y(N11121) );
  INVX1 gate3388 ( .A(N11062), .Y(N11122) );
  NAND2X1 gate3389 ( .A(N11062), .B(N9466), .Y(N11123) );
  NAND2X1 gate3390 ( .A(N11095), .B(N11066), .Y(N11124) );
  NAND2X1 gate3391 ( .A(N11098), .B(N11074), .Y(N11127) );
  NAND2X1 gate3392 ( .A(N11099), .B(N11076), .Y(N11130) );
  NAND2X1 gate3393 ( .A(N8687), .B(N11106), .Y(N11137) );
  NAND2X1 gate3394 ( .A(N8699), .B(N11108), .Y(N11138) );
  NAND2X1 gate3395 ( .A(N8766), .B(N11110), .Y(N11139) );
  NAND2X1 gate3396 ( .A(N8778), .B(N11112), .Y(N11140) );
  NAND2X1 gate3397 ( .A(N7456), .B(N11114), .Y(N11141) );
  NAND2X1 gate3398 ( .A(N7474), .B(N11116), .Y(N11142) );
  NAND2X1 gate3399 ( .A(N7512), .B(N11118), .Y(N11143) );
  NAND2X1 gate3400 ( .A(N7530), .B(N11120), .Y(N11144) );
  NAND2X1 gate3401 ( .A(N8705), .B(N11122), .Y(N11145) );
  AND2X1 gate3402_1 ( .A(N11103), .B(N8871), .Y(N11152_1) );
  AND2X1 gate3402 ( .A(N10283), .B(N11152_1), .Y(N11152) );
  AND2X1 gate3403_1 ( .A(N11100), .B(N7655), .Y(N11153_1) );
  AND2X1 gate3403 ( .A(N10283), .B(N11153_1), .Y(N11153) );
  AND2X1 gate3404_1 ( .A(N11103), .B(N9551), .Y(N11154_1) );
  AND2X1 gate3404 ( .A(N10119), .B(N11154_1), .Y(N11154) );
  AND2X1 gate3405_1 ( .A(N11100), .B(N9917), .Y(N11155_1) );
  AND2X1 gate3405 ( .A(N10119), .B(N11155_1), .Y(N11155) );
  NAND2X1 gate3406 ( .A(N11137), .B(N11107), .Y(N11156) );
  NAND2X1 gate3407 ( .A(N11138), .B(N11109), .Y(N11159) );
  NAND2X1 gate3408 ( .A(N11139), .B(N11111), .Y(N11162) );
  NAND2X1 gate3409 ( .A(N11140), .B(N11113), .Y(N11165) );
  NAND2X1 gate3410 ( .A(N11141), .B(N11115), .Y(N11168) );
  NAND2X1 gate3411 ( .A(N11142), .B(N11117), .Y(N11171) );
  NAND2X1 gate3412 ( .A(N11143), .B(N11119), .Y(N11174) );
  NAND2X1 gate3413 ( .A(N11144), .B(N11121), .Y(N11177) );
  NAND2X1 gate3414 ( .A(N11145), .B(N11123), .Y(N11180) );
  INVX1 gate3415 ( .A(N11124), .Y(N11183) );
  NAND2X1 gate3416 ( .A(N11124), .B(N9468), .Y(N11184) );
  INVX1 gate3417 ( .A(N11127), .Y(N11185) );
  NAND2X1 gate3418 ( .A(N11127), .B(N9508), .Y(N11186) );
  INVX1 gate3419 ( .A(N11130), .Y(N11187) );
  NAND2X1 gate3420 ( .A(N11130), .B(N9509), .Y(N11188) );
  OR2X1 gate3421_1 ( .A(N11152), .B(N11153), .Y(N11205_1) );
  OR2X1 gate3421_2 ( .A(N11154), .B(N11155), .Y(N11205_2) );
  OR2X1 gate3421 ( .A(N11205_1), .B(N11205_2), .Y(N11205) );
  NAND2X1 gate3422 ( .A(N8724), .B(N11183), .Y(N11210) );
  NAND2X1 gate3423 ( .A(N8790), .B(N11185), .Y(N11211) );
  NAND2X1 gate3424 ( .A(N8808), .B(N11187), .Y(N11212) );
  INVX1 gate3425 ( .A(N11168), .Y(N11213) );
  NAND2X1 gate3426 ( .A(N11168), .B(N8260), .Y(N11214) );
  INVX1 gate3427 ( .A(N11171), .Y(N11215) );
  NAND2X1 gate3428 ( .A(N11171), .B(N8261), .Y(N11216) );
  INVX1 gate3429 ( .A(N11174), .Y(N11217) );
  NAND2X1 gate3430 ( .A(N11174), .B(N8296), .Y(N11218) );
  INVX1 gate3431 ( .A(N11177), .Y(N11219) );
  NAND2X1 gate3432 ( .A(N11177), .B(N8297), .Y(N11220) );
  AND2X1 gate3433_1 ( .A(N11159), .B(N9575), .Y(N11222_1) );
  AND2X1 gate3433 ( .A(N1218), .B(N11222_1), .Y(N11222) );
  AND2X1 gate3434_1 ( .A(N11156), .B(N8927), .Y(N11223_1) );
  AND2X1 gate3434 ( .A(N1218), .B(N11223_1), .Y(N11223) );
  AND2X1 gate3435_1 ( .A(N11159), .B(N9935), .Y(N11224_1) );
  AND2X1 gate3435 ( .A(N750), .B(N11224_1), .Y(N11224) );
  AND2X1 gate3436_1 ( .A(N11156), .B(N10132), .Y(N11225_1) );
  AND2X1 gate3436 ( .A(N750), .B(N11225_1), .Y(N11225) );
  AND2X1 gate3437_1 ( .A(N11165), .B(N9608), .Y(N11226_1) );
  AND2X1 gate3437 ( .A(N10497), .B(N11226_1), .Y(N11226) );
  AND2X1 gate3438_1 ( .A(N11162), .B(N9001), .Y(N11227_1) );
  AND2X1 gate3438 ( .A(N10497), .B(N11227_1), .Y(N11227) );
  AND2X1 gate3439_1 ( .A(N11165), .B(N9949), .Y(N11228_1) );
  AND2X1 gate3439 ( .A(N10301), .B(N11228_1), .Y(N11228) );
  AND2X1 gate3440_1 ( .A(N11162), .B(N10160), .Y(N11229_1) );
  AND2X1 gate3440 ( .A(N10301), .B(N11229_1), .Y(N11229) );
  INVX1 gate3441 ( .A(N11180), .Y(N11231) );
  NAND2X1 gate3442 ( .A(N11180), .B(N9467), .Y(N11232) );
  NAND2X1 gate3443 ( .A(N11210), .B(N11184), .Y(N11233) );
  NAND2X1 gate3444 ( .A(N11211), .B(N11186), .Y(N11236) );
  NAND2X1 gate3445 ( .A(N11212), .B(N11188), .Y(N11239) );
  NAND2X1 gate3446 ( .A(N7459), .B(N11213), .Y(N11242) );
  NAND2X1 gate3447 ( .A(N7462), .B(N11215), .Y(N11243) );
  NAND2X1 gate3448 ( .A(N7515), .B(N11217), .Y(N11244) );
  NAND2X1 gate3449 ( .A(N7518), .B(N11219), .Y(N11245) );
  INVX1 gate3450 ( .A(N11205), .Y(N11246) );
  NAND2X1 gate3451 ( .A(N8708), .B(N11231), .Y(N11250) );
  OR2X1 gate3452_1 ( .A(N11222), .B(N11223), .Y(N11252_1) );
  OR2X1 gate3452_2 ( .A(N11224), .B(N11225), .Y(N11252_2) );
  OR2X1 gate3452 ( .A(N11252_1), .B(N11252_2), .Y(N11252) );
  OR2X1 gate3453_1 ( .A(N11226), .B(N11227), .Y(N11257_1) );
  OR2X1 gate3453_2 ( .A(N11228), .B(N11229), .Y(N11257_2) );
  OR2X1 gate3453 ( .A(N11257_1), .B(N11257_2), .Y(N11257) );
  NAND2X1 gate3454 ( .A(N11242), .B(N11214), .Y(N11260) );
  NAND2X1 gate3455 ( .A(N11243), .B(N11216), .Y(N11261) );
  NAND2X1 gate3456 ( .A(N11244), .B(N11218), .Y(N11262) );
  NAND2X1 gate3457 ( .A(N11245), .B(N11220), .Y(N11263) );
  INVX1 gate3458 ( .A(N11233), .Y(N11264) );
  NAND2X1 gate3459 ( .A(N11233), .B(N9322), .Y(N11265) );
  INVX1 gate3460 ( .A(N11236), .Y(N11267) );
  NAND2X1 gate3461 ( .A(N11236), .B(N9383), .Y(N11268) );
  INVX1 gate3462 ( .A(N11239), .Y(N11269) );
  NAND2X1 gate3463 ( .A(N11239), .B(N9384), .Y(N11270) );
  NAND2X1 gate3464 ( .A(N11250), .B(N11232), .Y(N11272) );
  INVX1 gate3465 ( .A(N11261), .Y(N11277) );
  AND2X1 gate3466 ( .A(N10273), .B(N11260), .Y(N11278) );
  INVX1 gate3467 ( .A(N11263), .Y(N11279) );
  AND2X1 gate3468 ( .A(N10119), .B(N11262), .Y(N11280) );
  NAND2X1 gate3469 ( .A(N8714), .B(N11264), .Y(N11282) );
  INVX1 gate3470 ( .A(N11252), .Y(N11283) );
  NAND2X1 gate3471 ( .A(N8793), .B(N11267), .Y(N11284) );
  NAND2X1 gate3472 ( .A(N8796), .B(N11269), .Y(N11285) );
  INVX1 gate3473 ( .A(N11257), .Y(N11286) );
  AND2X1 gate3474 ( .A(N11277), .B(N10479), .Y(N11288) );
  AND2X1 gate3475 ( .A(N11279), .B(N10283), .Y(N11289) );
  INVX1 gate3476 ( .A(N11272), .Y(N11290) );
  NAND2X1 gate3477 ( .A(N11272), .B(N9321), .Y(N11291) );
  NAND2X1 gate3478 ( .A(N11282), .B(N11265), .Y(N11292) );
  NAND2X1 gate3479 ( .A(N11284), .B(N11268), .Y(N11293) );
  NAND2X1 gate3480 ( .A(N11285), .B(N11270), .Y(N11294) );
  NAND2X1 gate3481 ( .A(N8711), .B(N11290), .Y(N11295) );
  INVX1 gate3482 ( .A(N11292), .Y(N11296) );
  INVX1 gate3483 ( .A(N11294), .Y(N11297) );
  AND2X1 gate3484 ( .A(N10301), .B(N11293), .Y(N11298) );
  OR2X1 gate3485 ( .A(N11288), .B(N11278), .Y(N11299) );
  OR2X1 gate3486 ( .A(N11289), .B(N11280), .Y(N11302) );
  NAND2X1 gate3487 ( .A(N11295), .B(N11291), .Y(N11307) );
  AND2X1 gate3488 ( .A(N11296), .B(N1218), .Y(N11308) );
  AND2X1 gate3489 ( .A(N11297), .B(N10497), .Y(N11309) );
  NAND2X1 gate3490 ( .A(N11302), .B(N11246), .Y(N11312) );
  NAND2X1 gate3491 ( .A(N11299), .B(N10836), .Y(N11313) );
  INVX1 gate3492 ( .A(N11299), .Y(N11314) );
  INVX1 gate3493 ( .A(N11302), .Y(N11315) );
  AND2X1 gate3494 ( .A(N750), .B(N11307), .Y(N11316) );
  OR2X1 gate3495 ( .A(N11309), .B(N11298), .Y(N11317) );
  NAND2X1 gate3496 ( .A(N11205), .B(N11315), .Y(N11320) );
  NAND2X1 gate3497 ( .A(N10739), .B(N11314), .Y(N11321) );
  OR2X1 gate3498 ( .A(N11308), .B(N11316), .Y(N11323) );
  NAND2X1 gate3499 ( .A(N11312), .B(N11320), .Y(N11327) );
  NAND2X1 gate3500 ( .A(N11313), .B(N11321), .Y(N11328) );
  NAND2X1 gate3501 ( .A(N11317), .B(N11286), .Y(N11329) );
  INVX1 gate3502 ( .A(N11317), .Y(N11331) );
  INVX1 gate3503 ( .A(N11327), .Y(N11333) );
  INVX1 gate3504 ( .A(N11328), .Y(N11334) );
  NAND2X1 gate3505 ( .A(N11257), .B(N11331), .Y(N11335) );
  NAND2X1 gate3506 ( .A(N11323), .B(N11283), .Y(N11336) );
  INVX1 gate3507 ( .A(N11323), .Y(N11337) );
  NAND2X1 gate3508 ( .A(N11329), .B(N11335), .Y(N11338) );
  NAND2X1 gate3509 ( .A(N11252), .B(N11337), .Y(N11339) );
  INVX1 gate3510 ( .A(N11338), .Y(N11340) );
  NAND2X1 gate3511 ( .A(N11336), .B(N11339), .Y(N11341) );
  INVX1 gate3512 ( .A(N11341), .Y(N11342) );
  BUFX2 gate3513 ( .A(N241_I), .Y(N241_O) );
endmodule



module c1908_synth ( N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, 
        N37, N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, 
        N82, N85, N88, N91, N94, N99, N104, N2753, N2754, N2755, N2756, N2762, 
        N2767, N2768, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, 
        N2787, N2811, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2899
 );
  input N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, N40, N43,
         N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, N85, N88,
         N91, N94, N99, N104;
  output N2753, N2754, N2755, N2756, N2762, N2767, N2768, N2779, N2780, N2781,
         N2782, N2783, N2784, N2785, N2786, N2787, N2811, N2886, N2887, N2888,
         N2889, N2890, N2891, N2892, N2899;
  wire   N190, N194, N197, N201, N206, N209, N212, N216, N220, N225, N229,
         N232, N235, N239, N243, N247, N251, N252, N253, N256, N257, N260,
         N263, N266, N269, N272, N275, N276, N277, N280, N283, N290, N297,
         N300, N303, N306, N313, N316, N319, N326, N331, N338, N343, N346,
         N349, N352, N355, N358, N361, N364, N367, N370, N373, N376, N379,
         N382, N385, N388, N534, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N559, N562, N565, N568, N571, N574, N577,
         N580, N583, N586, N589, N592, N595, N598, N601, N602, N603, N608,
         N612, N616, N619, N622, N625, N628, N631, N634, N637, N640, N643,
         N646, N649, N652, N655, N658, N661, N664, N667, N670, N673, N676,
         N679, N682, N685, N688, N691, N694, N697, N700, N703, N706, N709,
         N712, N715, N718, N721, N724, N727, N730, N733, N736, N739, N742,
         N745, N748, N751, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N903, N907, N910, N913, N914,
         N915, N916, N917, N918, N919, N920, N921, N922, N923, N926, N935,
         N938, N939, N942, N943, N946, N947, N950, N951, N954, N955, N958,
         N959, N962, N965, N968, N969, N972, N973, N976, N977, N980, N981,
         N984, N985, N988, N989, N990, N991, N992, N993, N994, N997, N998,
         N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010,
         N1013, N1016, N1019, N1022, N1025, N1028, N1031, N1034, N1037, N1040,
         N1043, N1046, N1049, N1054, N1055, N1063, N1064, N1067, N1068, N1119,
         N1120, N1121, N1122, N1128, N1129, N1130, N1131, N1132, N1133, N1148,
         N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158,
         N1159, N1160, N1161, N1162, N1163, N1164, N1167, N1168, N1171, N1188,
         N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214,
         N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224,
         N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1235, N1238,
         N1239, N1240, N1241, N1242, N1243, N1246, N1249, N1252, N1255, N1258,
         N1261, N1264, N1267, N1309, N1310, N1311, N1312, N1313, N1314, N1315,
         N1316, N1317, N1318, N1319, N1322, N1327, N1328, N1334, N1344, N1345,
         N1346, N1348, N1349, N1350, N1351, N1352, N1355, N1358, N1361, N1364,
         N1367, N1370, N1373, N1376, N1379, N1383, N1386, N1387, N1388, N1389,
         N1390, N1393, N1396, N1397, N1398, N1399, N1409, N1412, N1413, N1416,
         N1419, N1433, N1434, N1438, N1439, N1440, N1443, N1444, N1445, N1446,
         N1447, N1448, N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458,
         N1459, N1460, N1461, N1462, N1463, N1464, N1468, N1469, N1470, N1471,
         N1472, N1475, N1476, N1478, N1481, N1484, N1487, N1488, N1489, N1490,
         N1491, N1492, N1493, N1494, N1495, N1496, N1498, N1499, N1500, N1501,
         N1504, N1510, N1513, N1514, N1517, N1520, N1521, N1522, N1526, N1527,
         N1528, N1529, N1530, N1531, N1532, N1534, N1537, N1540, N1546, N1554,
         N1557, N1561, N1567, N1568, N1569, N1571, N1576, N1588, N1591, N1593,
         N1594, N1595, N1596, N1600, N1603, N1606, N1609, N1612, N1615, N1620,
         N1623, N1635, N1636, N1638, N1639, N1640, N1643, N1647, N1651, N1658,
         N1661, N1664, N1671, N1672, N1675, N1677, N1678, N1679, N1680, N1681,
         N1682, N1683, N1685, N1688, N1697, N1701, N1706, N1707, N1708, N1709,
         N1710, N1711, N1712, N1713, N1714, N1717, N1720, N1721, N1723, N1727,
         N1728, N1730, N1731, N1734, N1740, N1741, N1742, N1746, N1747, N1748,
         N1751, N1759, N1761, N1762, N1763, N1764, N1768, N1769, N1772, N1773,
         N1774, N1777, N1783, N1784, N1785, N1786, N1787, N1788, N1791, N1792,
         N1795, N1796, N1798, N1801, N1802, N1807, N1808, N1809, N1810, N1812,
         N1815, N1818, N1821, N1822, N1823, N1824, N1825, N1826, N1827, N1830,
         N1837, N1838, N1841, N1848, N1849, N1850, N1852, N1855, N1856, N1857,
         N1858, N1864, N1865, N1866, N1869, N1872, N1875, N1878, N1879, N1882,
         N1883, N1884, N1885, N1889, N1895, N1896, N1897, N1898, N1902, N1910,
         N1911, N1912, N1913, N1915, N1919, N1920, N1921, N1922, N1923, N1924,
         N1927, N1930, N1933, N1936, N1937, N1938, N1941, N1942, N1944, N1947,
         N1950, N1953, N1958, N1961, N1965, N1968, N1975, N1976, N1977, N1978,
         N1979, N1980, N1985, N1987, N1999, N2000, N2002, N2003, N2004, N2005,
         N2006, N2007, N2008, N2009, N2012, N2013, N2014, N2015, N2016, N2018,
         N2019, N2020, N2021, N2022, N2023, N2024, N2025, N2026, N2027, N2030,
         N2033, N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2047, N2052,
         N2055, N2060, N2061, N2062, N2067, N2068, N2071, N2076, N2077, N2078,
         N2081, N2086, N2089, N2104, N2119, N2129, N2143, N2148, N2151, N2196,
         N2199, N2202, N2205, N2214, N2215, N2216, N2217, N2222, N2223, N2224,
         N2225, N2226, N2227, N2228, N2229, N2230, N2231, N2232, N2233, N2234,
         N2235, N2236, N2237, N2240, N2241, N2244, N2245, N2250, N2253, N2256,
         N2257, N2260, N2263, N2266, N2269, N2272, N2279, N2286, N2297, N2315,
         N2326, N2340, N2353, N2361, N2375, N2384, N2385, N2386, N2426, N2427,
         N2537, N2540, N2543, N2546, N2549, N2552, N2555, N2558, N2561, N2564,
         N2567, N2570, N2573, N2576, N2594, N2597, N2600, N2603, N2606, N2611,
         N2614, N2617, N2620, N2627, N2628, N2629, N2630, N2631, N2632, N2633,
         N2634, N2639, N2642, N2645, N2648, N2651, N2655, N2658, N2661, N2664,
         N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2682, N2683,
         N2688, N2689, N2690, N2691, N2710, N2720, N2721, N2722, N2723, N2724,
         N2725, N2726, N2727, N2728, N2729, N2730, N2731, N2732, N2733, N2734,
         N2735, N2736, N2737, N2738, N2739, N2740, N2741, N2742, N2743, N2744,
         N2745, N2746, N2747, N2750, N2757, N2758, N2759, N2760, N2761, N2763,
         N2764, N2765, N2766, N2773, N2776, N2788, N2789, N2800, N2807, N2808,
         N2809, N2810, N2812, N2815, N2818, N2821, N2824, N2827, N2828, N2829,
         N2843, N2846, N2850, N2851, N2852, N2853, N2854, N2857, N2858, N2859,
         N2860, N2861, N2862, N2863, N2866, N2867, N2868, N2869, N2870, N2871,
         N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880, N2881,
         N2882, N2883, N2895, N2896, N2897, N2898, N592_1, N643_1, N655_1,
         N724_1, N921_1, N921_2, N922_1, N922_2, N926_1, N2279_1, N2279_2,
         N2279_3, N2384_1, N2384_2, N2537_1, N2537_2, N2540_1, N2540_2,
         N2543_1, N2543_2, N2546_1, N2546_2, N2549_1, N2549_2, N2552_1,
         N2552_2, N2555_1, N2555_2, N2558_1, N2558_2, N2558_3, N2561_1,
         N2561_2, N2561_3, N2564_1, N2564_2, N2564_3, N2567_1, N2567_2,
         N2567_3, N2570_1, N2570_2, N2570_3, N2573_1, N2573_2, N2573_3,
         N2576_1, N2576_2, N2576_3, N2594_1, N2594_2, N2597_1, N2597_2,
         N2600_1, N2600_2, N2603_1, N2603_2, N2606_1, N2606_2, N2611_1,
         N2611_2, N2614_1, N2614_2, N2617_1, N2617_2, N2620_1, N2620_2,
         N2627_1, N2627_2, N2628_1, N2628_2, N2629_1, N2629_2, N2630_1,
         N2630_2, N2631_1, N2631_2, N2632_1, N2632_2, N2633_1, N2633_2,
         N2634_1, N2634_2, N2639_1, N2639_2, N2639_3, N2642_1, N2642_2,
         N2642_3, N2645_1, N2645_2, N2645_3, N2648_1, N2648_2, N2648_3,
         N2651_1, N2651_2, N2651_3, N2655_1, N2655_2, N2655_3, N2658_1,
         N2658_2, N2658_3, N2661_1, N2661_2, N2661_3, N2664_1, N2664_2,
         N2664_3, N2710_1, N2710_2, N2710_3, N2710_4, N2710_5, N2710_6,
         N2745_1, N2745_2, N2745_3, N2746_1, N2746_2, N2746_3, N2747_1,
         N2747_2, N2747_3, N2747_4, N2747_5, N2747_6, N2750_1, N2750_2,
         N2750_3, N2750_4, N2750_5, N2750_6, N2788_1, N2800_1, N2800_2,
         N2812_1, N2815_1, N2818_1, N2821_1, N2824_1, N2829_1;

  INVX1 gate1 ( .A(N1), .Y(N190) );
  INVX1 gate2 ( .A(N4), .Y(N194) );
  INVX1 gate3 ( .A(N7), .Y(N197) );
  INVX1 gate4 ( .A(N10), .Y(N201) );
  INVX1 gate5 ( .A(N13), .Y(N206) );
  INVX1 gate6 ( .A(N16), .Y(N209) );
  INVX1 gate7 ( .A(N19), .Y(N212) );
  INVX1 gate8 ( .A(N22), .Y(N216) );
  INVX1 gate9 ( .A(N25), .Y(N220) );
  INVX1 gate10 ( .A(N28), .Y(N225) );
  INVX1 gate11 ( .A(N31), .Y(N229) );
  INVX1 gate12 ( .A(N34), .Y(N232) );
  INVX1 gate13 ( .A(N37), .Y(N235) );
  INVX1 gate14 ( .A(N40), .Y(N239) );
  INVX1 gate15 ( .A(N43), .Y(N243) );
  INVX1 gate16 ( .A(N46), .Y(N247) );
  NAND2X1 gate17 ( .A(N63), .B(N88), .Y(N251) );
  NAND2X1 gate18 ( .A(N66), .B(N91), .Y(N252) );
  INVX1 gate19 ( .A(N72), .Y(N253) );
  INVX1 gate20 ( .A(N72), .Y(N256) );
  BUFX2 gate21 ( .A(N69), .Y(N257) );
  BUFX2 gate22 ( .A(N69), .Y(N260) );
  INVX1 gate23 ( .A(N76), .Y(N263) );
  INVX1 gate24 ( .A(N79), .Y(N266) );
  INVX1 gate25 ( .A(N82), .Y(N269) );
  INVX1 gate26 ( .A(N85), .Y(N272) );
  INVX1 gate27 ( .A(N104), .Y(N275) );
  INVX1 gate28 ( .A(N104), .Y(N276) );
  INVX1 gate29 ( .A(N88), .Y(N277) );
  INVX1 gate30 ( .A(N91), .Y(N280) );
  BUFX2 gate31 ( .A(N94), .Y(N283) );
  INVX1 gate32 ( .A(N94), .Y(N290) );
  BUFX2 gate33 ( .A(N94), .Y(N297) );
  INVX1 gate34 ( .A(N94), .Y(N300) );
  BUFX2 gate35 ( .A(N99), .Y(N303) );
  INVX1 gate36 ( .A(N99), .Y(N306) );
  INVX1 gate37 ( .A(N99), .Y(N313) );
  BUFX2 gate38 ( .A(N104), .Y(N316) );
  INVX1 gate39 ( .A(N104), .Y(N319) );
  BUFX2 gate40 ( .A(N104), .Y(N326) );
  BUFX2 gate41 ( .A(N104), .Y(N331) );
  INVX1 gate42 ( .A(N104), .Y(N338) );
  BUFX2 gate43 ( .A(N1), .Y(N343) );
  BUFX2 gate44 ( .A(N4), .Y(N346) );
  BUFX2 gate45 ( .A(N7), .Y(N349) );
  BUFX2 gate46 ( .A(N10), .Y(N352) );
  BUFX2 gate47 ( .A(N13), .Y(N355) );
  BUFX2 gate48 ( .A(N16), .Y(N358) );
  BUFX2 gate49 ( .A(N19), .Y(N361) );
  BUFX2 gate50 ( .A(N22), .Y(N364) );
  BUFX2 gate51 ( .A(N25), .Y(N367) );
  BUFX2 gate52 ( .A(N28), .Y(N370) );
  BUFX2 gate53 ( .A(N31), .Y(N373) );
  BUFX2 gate54 ( .A(N34), .Y(N376) );
  BUFX2 gate55 ( .A(N37), .Y(N379) );
  BUFX2 gate56 ( .A(N40), .Y(N382) );
  BUFX2 gate57 ( .A(N43), .Y(N385) );
  BUFX2 gate58 ( .A(N46), .Y(N388) );
  INVX1 gate59 ( .A(N343), .Y(N534) );
  INVX1 gate60 ( .A(N346), .Y(N535) );
  INVX1 gate61 ( .A(N349), .Y(N536) );
  INVX1 gate62 ( .A(N352), .Y(N537) );
  INVX1 gate63 ( .A(N355), .Y(N538) );
  INVX1 gate64 ( .A(N358), .Y(N539) );
  INVX1 gate65 ( .A(N361), .Y(N540) );
  INVX1 gate66 ( .A(N364), .Y(N541) );
  INVX1 gate67 ( .A(N367), .Y(N542) );
  INVX1 gate68 ( .A(N370), .Y(N543) );
  INVX1 gate69 ( .A(N373), .Y(N544) );
  INVX1 gate70 ( .A(N376), .Y(N545) );
  INVX1 gate71 ( .A(N379), .Y(N546) );
  INVX1 gate72 ( .A(N382), .Y(N547) );
  INVX1 gate73 ( .A(N385), .Y(N548) );
  INVX1 gate74 ( .A(N388), .Y(N549) );
  NAND2X1 gate75 ( .A(N306), .B(N331), .Y(N550) );
  NAND2X1 gate76 ( .A(N306), .B(N331), .Y(N551) );
  NAND2X1 gate77 ( .A(N306), .B(N331), .Y(N552) );
  NAND2X1 gate78 ( .A(N306), .B(N331), .Y(N553) );
  NAND2X1 gate79 ( .A(N306), .B(N331), .Y(N554) );
  NAND2X1 gate80 ( .A(N306), .B(N331), .Y(N555) );
  BUFX2 gate81 ( .A(N190), .Y(N556) );
  BUFX2 gate82 ( .A(N194), .Y(N559) );
  BUFX2 gate83 ( .A(N206), .Y(N562) );
  BUFX2 gate84 ( .A(N209), .Y(N565) );
  BUFX2 gate85 ( .A(N225), .Y(N568) );
  BUFX2 gate86 ( .A(N243), .Y(N571) );
  AND2X1 gate87 ( .A(N63), .B(N319), .Y(N574) );
  BUFX2 gate88 ( .A(N220), .Y(N577) );
  BUFX2 gate89 ( .A(N229), .Y(N580) );
  BUFX2 gate90 ( .A(N232), .Y(N583) );
  AND2X1 gate91 ( .A(N66), .B(N319), .Y(N586) );
  BUFX2 gate92 ( .A(N239), .Y(N589) );
  AND2X1 gate93_1 ( .A(N49), .B(N253), .Y(N592_1) );
  AND2X1 gate93 ( .A(N319), .B(N592_1), .Y(N592) );
  BUFX2 gate94 ( .A(N247), .Y(N595) );
  BUFX2 gate95 ( .A(N239), .Y(N598) );
  NAND2X1 gate96 ( .A(N326), .B(N277), .Y(N601) );
  NAND2X1 gate97 ( .A(N326), .B(N280), .Y(N602) );
  NAND2X1 gate98 ( .A(N260), .B(N72), .Y(N603) );
  NAND2X1 gate99 ( .A(N260), .B(N300), .Y(N608) );
  NAND2X1 gate100 ( .A(N256), .B(N300), .Y(N612) );
  BUFX2 gate101 ( .A(N201), .Y(N616) );
  BUFX2 gate102 ( .A(N216), .Y(N619) );
  BUFX2 gate103 ( .A(N220), .Y(N622) );
  BUFX2 gate104 ( .A(N239), .Y(N625) );
  BUFX2 gate105 ( .A(N190), .Y(N628) );
  BUFX2 gate106 ( .A(N190), .Y(N631) );
  BUFX2 gate107 ( .A(N194), .Y(N634) );
  BUFX2 gate108 ( .A(N229), .Y(N637) );
  BUFX2 gate109 ( .A(N197), .Y(N640) );
  AND2X1 gate110_1 ( .A(N56), .B(N257), .Y(N643_1) );
  AND2X1 gate110 ( .A(N319), .B(N643_1), .Y(N643) );
  BUFX2 gate111 ( .A(N232), .Y(N646) );
  BUFX2 gate112 ( .A(N201), .Y(N649) );
  BUFX2 gate113 ( .A(N235), .Y(N652) );
  AND2X1 gate114_1 ( .A(N60), .B(N257), .Y(N655_1) );
  AND2X1 gate114 ( .A(N319), .B(N655_1), .Y(N655) );
  BUFX2 gate115 ( .A(N263), .Y(N658) );
  BUFX2 gate116 ( .A(N263), .Y(N661) );
  BUFX2 gate117 ( .A(N266), .Y(N664) );
  BUFX2 gate118 ( .A(N266), .Y(N667) );
  BUFX2 gate119 ( .A(N269), .Y(N670) );
  BUFX2 gate120 ( .A(N269), .Y(N673) );
  BUFX2 gate121 ( .A(N272), .Y(N676) );
  BUFX2 gate122 ( .A(N272), .Y(N679) );
  AND2X1 gate123 ( .A(N251), .B(N316), .Y(N682) );
  AND2X1 gate124 ( .A(N252), .B(N316), .Y(N685) );
  BUFX2 gate125 ( .A(N197), .Y(N688) );
  BUFX2 gate126 ( .A(N197), .Y(N691) );
  BUFX2 gate127 ( .A(N212), .Y(N694) );
  BUFX2 gate128 ( .A(N212), .Y(N697) );
  BUFX2 gate129 ( .A(N247), .Y(N700) );
  BUFX2 gate130 ( .A(N247), .Y(N703) );
  BUFX2 gate131 ( .A(N235), .Y(N706) );
  BUFX2 gate132 ( .A(N235), .Y(N709) );
  BUFX2 gate133 ( .A(N201), .Y(N712) );
  BUFX2 gate134 ( .A(N201), .Y(N715) );
  BUFX2 gate135 ( .A(N206), .Y(N718) );
  BUFX2 gate136 ( .A(N216), .Y(N721) );
  AND2X1 gate137_1 ( .A(N53), .B(N253), .Y(N724_1) );
  AND2X1 gate137 ( .A(N319), .B(N724_1), .Y(N724) );
  BUFX2 gate138 ( .A(N243), .Y(N727) );
  BUFX2 gate139 ( .A(N220), .Y(N730) );
  BUFX2 gate140 ( .A(N220), .Y(N733) );
  BUFX2 gate141 ( .A(N209), .Y(N736) );
  BUFX2 gate142 ( .A(N216), .Y(N739) );
  BUFX2 gate143 ( .A(N225), .Y(N742) );
  BUFX2 gate144 ( .A(N243), .Y(N745) );
  BUFX2 gate145 ( .A(N212), .Y(N748) );
  BUFX2 gate146 ( .A(N225), .Y(N751) );
  INVX1 gate147 ( .A(N682), .Y(N886) );
  INVX1 gate148 ( .A(N685), .Y(N887) );
  INVX1 gate149 ( .A(N616), .Y(N888) );
  INVX1 gate150 ( .A(N619), .Y(N889) );
  INVX1 gate151 ( .A(N622), .Y(N890) );
  INVX1 gate152 ( .A(N625), .Y(N891) );
  INVX1 gate153 ( .A(N631), .Y(N892) );
  INVX1 gate154 ( .A(N643), .Y(N893) );
  INVX1 gate155 ( .A(N649), .Y(N894) );
  INVX1 gate156 ( .A(N652), .Y(N895) );
  INVX1 gate157 ( .A(N655), .Y(N896) );
  AND2X1 gate158 ( .A(N49), .B(N612), .Y(N897) );
  AND2X1 gate159 ( .A(N56), .B(N608), .Y(N898) );
  NAND2X1 gate160 ( .A(N53), .B(N612), .Y(N899) );
  NAND2X1 gate161 ( .A(N60), .B(N608), .Y(N903) );
  NAND2X1 gate162 ( .A(N49), .B(N612), .Y(N907) );
  NAND2X1 gate163 ( .A(N56), .B(N608), .Y(N910) );
  INVX1 gate164 ( .A(N661), .Y(N913) );
  INVX1 gate165 ( .A(N658), .Y(N914) );
  INVX1 gate166 ( .A(N667), .Y(N915) );
  INVX1 gate167 ( .A(N664), .Y(N916) );
  INVX1 gate168 ( .A(N673), .Y(N917) );
  INVX1 gate169 ( .A(N670), .Y(N918) );
  INVX1 gate170 ( .A(N679), .Y(N919) );
  INVX1 gate171 ( .A(N676), .Y(N920) );
  NAND2X1 gate172_1 ( .A(N277), .B(N297), .Y(N921_1) );
  NAND2X1 gate172_2 ( .A(N326), .B(N603), .Y(N921_2) );
  NAND2X1 gate172 ( .A(N921_1), .B(N921_2), .Y(N921) );
  NAND2X1 gate173_1 ( .A(N280), .B(N297), .Y(N922_1) );
  NAND2X1 gate173_2 ( .A(N326), .B(N603), .Y(N922_2) );
  NAND2X1 gate173 ( .A(N922_1), .B(N922_2), .Y(N922) );
  NAND3X1 gate174 ( .A(N303), .B(N338), .C(N603), .Y(N923) );
  AND2X1 gate175_1 ( .A(N303), .B(N338), .Y(N926_1) );
  AND2X1 gate175 ( .A(N603), .B(N926_1), .Y(N926) );
  BUFX2 gate176 ( .A(N556), .Y(N935) );
  INVX1 gate177 ( .A(N688), .Y(N938) );
  BUFX2 gate178 ( .A(N556), .Y(N939) );
  INVX1 gate179 ( .A(N691), .Y(N942) );
  BUFX2 gate180 ( .A(N562), .Y(N943) );
  INVX1 gate181 ( .A(N694), .Y(N946) );
  BUFX2 gate182 ( .A(N562), .Y(N947) );
  INVX1 gate183 ( .A(N697), .Y(N950) );
  BUFX2 gate184 ( .A(N568), .Y(N951) );
  INVX1 gate185 ( .A(N700), .Y(N954) );
  BUFX2 gate186 ( .A(N568), .Y(N955) );
  INVX1 gate187 ( .A(N703), .Y(N958) );
  BUFX2 gate188 ( .A(N574), .Y(N959) );
  BUFX2 gate189 ( .A(N574), .Y(N962) );
  BUFX2 gate190 ( .A(N580), .Y(N965) );
  INVX1 gate191 ( .A(N706), .Y(N968) );
  BUFX2 gate192 ( .A(N580), .Y(N969) );
  INVX1 gate193 ( .A(N709), .Y(N972) );
  BUFX2 gate194 ( .A(N586), .Y(N973) );
  INVX1 gate195 ( .A(N712), .Y(N976) );
  BUFX2 gate196 ( .A(N586), .Y(N977) );
  INVX1 gate197 ( .A(N715), .Y(N980) );
  BUFX2 gate198 ( .A(N592), .Y(N981) );
  INVX1 gate199 ( .A(N628), .Y(N984) );
  BUFX2 gate200 ( .A(N592), .Y(N985) );
  INVX1 gate201 ( .A(N718), .Y(N988) );
  INVX1 gate202 ( .A(N721), .Y(N989) );
  INVX1 gate203 ( .A(N634), .Y(N990) );
  INVX1 gate204 ( .A(N724), .Y(N991) );
  INVX1 gate205 ( .A(N727), .Y(N992) );
  INVX1 gate206 ( .A(N637), .Y(N993) );
  BUFX2 gate207 ( .A(N595), .Y(N994) );
  INVX1 gate208 ( .A(N730), .Y(N997) );
  BUFX2 gate209 ( .A(N595), .Y(N998) );
  INVX1 gate210 ( .A(N733), .Y(N1001) );
  INVX1 gate211 ( .A(N736), .Y(N1002) );
  INVX1 gate212 ( .A(N739), .Y(N1003) );
  INVX1 gate213 ( .A(N640), .Y(N1004) );
  INVX1 gate214 ( .A(N742), .Y(N1005) );
  INVX1 gate215 ( .A(N745), .Y(N1006) );
  INVX1 gate216 ( .A(N646), .Y(N1007) );
  INVX1 gate217 ( .A(N748), .Y(N1008) );
  INVX1 gate218 ( .A(N751), .Y(N1009) );
  BUFX2 gate219 ( .A(N559), .Y(N1010) );
  BUFX2 gate220 ( .A(N559), .Y(N1013) );
  BUFX2 gate221 ( .A(N565), .Y(N1016) );
  BUFX2 gate222 ( .A(N565), .Y(N1019) );
  BUFX2 gate223 ( .A(N571), .Y(N1022) );
  BUFX2 gate224 ( .A(N571), .Y(N1025) );
  BUFX2 gate225 ( .A(N577), .Y(N1028) );
  BUFX2 gate226 ( .A(N577), .Y(N1031) );
  BUFX2 gate227 ( .A(N583), .Y(N1034) );
  BUFX2 gate228 ( .A(N583), .Y(N1037) );
  BUFX2 gate229 ( .A(N589), .Y(N1040) );
  BUFX2 gate230 ( .A(N589), .Y(N1043) );
  BUFX2 gate231 ( .A(N598), .Y(N1046) );
  BUFX2 gate232 ( .A(N598), .Y(N1049) );
  NAND2X1 gate233 ( .A(N619), .B(N888), .Y(N1054) );
  NAND2X1 gate234 ( .A(N616), .B(N889), .Y(N1055) );
  NAND2X1 gate235 ( .A(N625), .B(N890), .Y(N1063) );
  NAND2X1 gate236 ( .A(N622), .B(N891), .Y(N1064) );
  NAND2X1 gate237 ( .A(N655), .B(N895), .Y(N1067) );
  NAND2X1 gate238 ( .A(N652), .B(N896), .Y(N1068) );
  NAND2X1 gate239 ( .A(N721), .B(N988), .Y(N1119) );
  NAND2X1 gate240 ( .A(N718), .B(N989), .Y(N1120) );
  NAND2X1 gate241 ( .A(N727), .B(N991), .Y(N1121) );
  NAND2X1 gate242 ( .A(N724), .B(N992), .Y(N1122) );
  NAND2X1 gate243 ( .A(N739), .B(N1002), .Y(N1128) );
  NAND2X1 gate244 ( .A(N736), .B(N1003), .Y(N1129) );
  NAND2X1 gate245 ( .A(N745), .B(N1005), .Y(N1130) );
  NAND2X1 gate246 ( .A(N742), .B(N1006), .Y(N1131) );
  NAND2X1 gate247 ( .A(N751), .B(N1008), .Y(N1132) );
  NAND2X1 gate248 ( .A(N748), .B(N1009), .Y(N1133) );
  INVX1 gate249 ( .A(N939), .Y(N1148) );
  INVX1 gate250 ( .A(N935), .Y(N1149) );
  NAND2X1 gate251 ( .A(N1054), .B(N1055), .Y(N1150) );
  INVX1 gate252 ( .A(N943), .Y(N1151) );
  INVX1 gate253 ( .A(N947), .Y(N1152) );
  INVX1 gate254 ( .A(N955), .Y(N1153) );
  INVX1 gate255 ( .A(N951), .Y(N1154) );
  INVX1 gate256 ( .A(N962), .Y(N1155) );
  INVX1 gate257 ( .A(N969), .Y(N1156) );
  INVX1 gate258 ( .A(N977), .Y(N1157) );
  NAND2X1 gate259 ( .A(N1063), .B(N1064), .Y(N1158) );
  INVX1 gate260 ( .A(N985), .Y(N1159) );
  NAND2X1 gate261 ( .A(N985), .B(N892), .Y(N1160) );
  INVX1 gate262 ( .A(N998), .Y(N1161) );
  NAND2X1 gate263 ( .A(N1067), .B(N1068), .Y(N1162) );
  INVX1 gate264 ( .A(N899), .Y(N1163) );
  BUFX2 gate265 ( .A(N899), .Y(N1164) );
  INVX1 gate266 ( .A(N903), .Y(N1167) );
  BUFX2 gate267 ( .A(N903), .Y(N1168) );
  NAND2X1 gate268 ( .A(N921), .B(N923), .Y(N1171) );
  NAND2X1 gate269 ( .A(N922), .B(N923), .Y(N1188) );
  INVX1 gate270 ( .A(N1010), .Y(N1205) );
  NAND2X1 gate271 ( .A(N1010), .B(N938), .Y(N1206) );
  INVX1 gate272 ( .A(N1013), .Y(N1207) );
  NAND2X1 gate273 ( .A(N1013), .B(N942), .Y(N1208) );
  INVX1 gate274 ( .A(N1016), .Y(N1209) );
  NAND2X1 gate275 ( .A(N1016), .B(N946), .Y(N1210) );
  INVX1 gate276 ( .A(N1019), .Y(N1211) );
  NAND2X1 gate277 ( .A(N1019), .B(N950), .Y(N1212) );
  INVX1 gate278 ( .A(N1022), .Y(N1213) );
  NAND2X1 gate279 ( .A(N1022), .B(N954), .Y(N1214) );
  INVX1 gate280 ( .A(N1025), .Y(N1215) );
  NAND2X1 gate281 ( .A(N1025), .B(N958), .Y(N1216) );
  INVX1 gate282 ( .A(N1028), .Y(N1217) );
  INVX1 gate283 ( .A(N959), .Y(N1218) );
  INVX1 gate284 ( .A(N1031), .Y(N1219) );
  INVX1 gate285 ( .A(N1034), .Y(N1220) );
  NAND2X1 gate286 ( .A(N1034), .B(N968), .Y(N1221) );
  INVX1 gate287 ( .A(N965), .Y(N1222) );
  INVX1 gate288 ( .A(N1037), .Y(N1223) );
  NAND2X1 gate289 ( .A(N1037), .B(N972), .Y(N1224) );
  INVX1 gate290 ( .A(N1040), .Y(N1225) );
  NAND2X1 gate291 ( .A(N1040), .B(N976), .Y(N1226) );
  INVX1 gate292 ( .A(N973), .Y(N1227) );
  INVX1 gate293 ( .A(N1043), .Y(N1228) );
  NAND2X1 gate294 ( .A(N1043), .B(N980), .Y(N1229) );
  INVX1 gate295 ( .A(N981), .Y(N1230) );
  NAND2X1 gate296 ( .A(N981), .B(N984), .Y(N1231) );
  NAND2X1 gate297 ( .A(N1119), .B(N1120), .Y(N1232) );
  NAND2X1 gate298 ( .A(N1121), .B(N1122), .Y(N1235) );
  INVX1 gate299 ( .A(N1046), .Y(N1238) );
  NAND2X1 gate300 ( .A(N1046), .B(N997), .Y(N1239) );
  INVX1 gate301 ( .A(N994), .Y(N1240) );
  INVX1 gate302 ( .A(N1049), .Y(N1241) );
  NAND2X1 gate303 ( .A(N1049), .B(N1001), .Y(N1242) );
  NAND2X1 gate304 ( .A(N1128), .B(N1129), .Y(N1243) );
  NAND2X1 gate305 ( .A(N1130), .B(N1131), .Y(N1246) );
  NAND2X1 gate306 ( .A(N1132), .B(N1133), .Y(N1249) );
  BUFX2 gate307 ( .A(N907), .Y(N1252) );
  BUFX2 gate308 ( .A(N907), .Y(N1255) );
  BUFX2 gate309 ( .A(N910), .Y(N1258) );
  BUFX2 gate310 ( .A(N910), .Y(N1261) );
  INVX1 gate311 ( .A(N1150), .Y(N1264) );
  NAND2X1 gate312 ( .A(N631), .B(N1159), .Y(N1267) );
  NAND2X1 gate313 ( .A(N688), .B(N1205), .Y(N1309) );
  NAND2X1 gate314 ( .A(N691), .B(N1207), .Y(N1310) );
  NAND2X1 gate315 ( .A(N694), .B(N1209), .Y(N1311) );
  NAND2X1 gate316 ( .A(N697), .B(N1211), .Y(N1312) );
  NAND2X1 gate317 ( .A(N700), .B(N1213), .Y(N1313) );
  NAND2X1 gate318 ( .A(N703), .B(N1215), .Y(N1314) );
  NAND2X1 gate319 ( .A(N706), .B(N1220), .Y(N1315) );
  NAND2X1 gate320 ( .A(N709), .B(N1223), .Y(N1316) );
  NAND2X1 gate321 ( .A(N712), .B(N1225), .Y(N1317) );
  NAND2X1 gate322 ( .A(N715), .B(N1228), .Y(N1318) );
  INVX1 gate323 ( .A(N1158), .Y(N1319) );
  NAND2X1 gate324 ( .A(N628), .B(N1230), .Y(N1322) );
  NAND2X1 gate325 ( .A(N730), .B(N1238), .Y(N1327) );
  NAND2X1 gate326 ( .A(N733), .B(N1241), .Y(N1328) );
  INVX1 gate327 ( .A(N1162), .Y(N1334) );
  NAND2X1 gate328 ( .A(N1267), .B(N1160), .Y(N1344) );
  NAND2X1 gate329 ( .A(N1249), .B(N894), .Y(N1345) );
  INVX1 gate330 ( .A(N1249), .Y(N1346) );
  INVX1 gate331 ( .A(N1255), .Y(N1348) );
  INVX1 gate332 ( .A(N1252), .Y(N1349) );
  INVX1 gate333 ( .A(N1261), .Y(N1350) );
  INVX1 gate334 ( .A(N1258), .Y(N1351) );
  NAND2X1 gate335 ( .A(N1309), .B(N1206), .Y(N1352) );
  NAND2X1 gate336 ( .A(N1310), .B(N1208), .Y(N1355) );
  NAND2X1 gate337 ( .A(N1311), .B(N1210), .Y(N1358) );
  NAND2X1 gate338 ( .A(N1312), .B(N1212), .Y(N1361) );
  NAND2X1 gate339 ( .A(N1313), .B(N1214), .Y(N1364) );
  NAND2X1 gate340 ( .A(N1314), .B(N1216), .Y(N1367) );
  NAND2X1 gate341 ( .A(N1315), .B(N1221), .Y(N1370) );
  NAND2X1 gate342 ( .A(N1316), .B(N1224), .Y(N1373) );
  NAND2X1 gate343 ( .A(N1317), .B(N1226), .Y(N1376) );
  NAND2X1 gate344 ( .A(N1318), .B(N1229), .Y(N1379) );
  NAND2X1 gate345 ( .A(N1322), .B(N1231), .Y(N1383) );
  INVX1 gate346 ( .A(N1232), .Y(N1386) );
  NAND2X1 gate347 ( .A(N1232), .B(N990), .Y(N1387) );
  INVX1 gate348 ( .A(N1235), .Y(N1388) );
  NAND2X1 gate349 ( .A(N1235), .B(N993), .Y(N1389) );
  NAND2X1 gate350 ( .A(N1327), .B(N1239), .Y(N1390) );
  NAND2X1 gate351 ( .A(N1328), .B(N1242), .Y(N1393) );
  INVX1 gate352 ( .A(N1243), .Y(N1396) );
  NAND2X1 gate353 ( .A(N1243), .B(N1004), .Y(N1397) );
  INVX1 gate354 ( .A(N1246), .Y(N1398) );
  NAND2X1 gate355 ( .A(N1246), .B(N1007), .Y(N1399) );
  INVX1 gate356 ( .A(N1319), .Y(N1409) );
  NAND2X1 gate357 ( .A(N649), .B(N1346), .Y(N1412) );
  INVX1 gate358 ( .A(N1334), .Y(N1413) );
  BUFX2 gate359 ( .A(N1264), .Y(N1416) );
  BUFX2 gate360 ( .A(N1264), .Y(N1419) );
  NAND2X1 gate361 ( .A(N634), .B(N1386), .Y(N1433) );
  NAND2X1 gate362 ( .A(N637), .B(N1388), .Y(N1434) );
  NAND2X1 gate363 ( .A(N640), .B(N1396), .Y(N1438) );
  NAND2X1 gate364 ( .A(N646), .B(N1398), .Y(N1439) );
  INVX1 gate365 ( .A(N1344), .Y(N1440) );
  NAND2X1 gate366 ( .A(N1355), .B(N1148), .Y(N1443) );
  INVX1 gate367 ( .A(N1355), .Y(N1444) );
  NAND2X1 gate368 ( .A(N1352), .B(N1149), .Y(N1445) );
  INVX1 gate369 ( .A(N1352), .Y(N1446) );
  NAND2X1 gate370 ( .A(N1358), .B(N1151), .Y(N1447) );
  INVX1 gate371 ( .A(N1358), .Y(N1448) );
  NAND2X1 gate372 ( .A(N1361), .B(N1152), .Y(N1451) );
  INVX1 gate373 ( .A(N1361), .Y(N1452) );
  NAND2X1 gate374 ( .A(N1367), .B(N1153), .Y(N1453) );
  INVX1 gate375 ( .A(N1367), .Y(N1454) );
  NAND2X1 gate376 ( .A(N1364), .B(N1154), .Y(N1455) );
  INVX1 gate377 ( .A(N1364), .Y(N1456) );
  NAND2X1 gate378 ( .A(N1373), .B(N1156), .Y(N1457) );
  INVX1 gate379 ( .A(N1373), .Y(N1458) );
  NAND2X1 gate380 ( .A(N1379), .B(N1157), .Y(N1459) );
  INVX1 gate381 ( .A(N1379), .Y(N1460) );
  INVX1 gate382 ( .A(N1383), .Y(N1461) );
  NAND2X1 gate383 ( .A(N1393), .B(N1161), .Y(N1462) );
  INVX1 gate384 ( .A(N1393), .Y(N1463) );
  NAND2X1 gate385 ( .A(N1345), .B(N1412), .Y(N1464) );
  INVX1 gate386 ( .A(N1370), .Y(N1468) );
  NAND2X1 gate387 ( .A(N1370), .B(N1222), .Y(N1469) );
  INVX1 gate388 ( .A(N1376), .Y(N1470) );
  NAND2X1 gate389 ( .A(N1376), .B(N1227), .Y(N1471) );
  NAND2X1 gate390 ( .A(N1387), .B(N1433), .Y(N1472) );
  INVX1 gate391 ( .A(N1390), .Y(N1475) );
  NAND2X1 gate392 ( .A(N1390), .B(N1240), .Y(N1476) );
  NAND2X1 gate393 ( .A(N1389), .B(N1434), .Y(N1478) );
  NAND2X1 gate394 ( .A(N1399), .B(N1439), .Y(N1481) );
  NAND2X1 gate395 ( .A(N1397), .B(N1438), .Y(N1484) );
  NAND2X1 gate396 ( .A(N939), .B(N1444), .Y(N1487) );
  NAND2X1 gate397 ( .A(N935), .B(N1446), .Y(N1488) );
  NAND2X1 gate398 ( .A(N943), .B(N1448), .Y(N1489) );
  INVX1 gate399 ( .A(N1419), .Y(N1490) );
  INVX1 gate400 ( .A(N1416), .Y(N1491) );
  NAND2X1 gate401 ( .A(N947), .B(N1452), .Y(N1492) );
  NAND2X1 gate402 ( .A(N955), .B(N1454), .Y(N1493) );
  NAND2X1 gate403 ( .A(N951), .B(N1456), .Y(N1494) );
  NAND2X1 gate404 ( .A(N969), .B(N1458), .Y(N1495) );
  NAND2X1 gate405 ( .A(N977), .B(N1460), .Y(N1496) );
  NAND2X1 gate406 ( .A(N998), .B(N1463), .Y(N1498) );
  INVX1 gate407 ( .A(N1440), .Y(N1499) );
  NAND2X1 gate408 ( .A(N965), .B(N1468), .Y(N1500) );
  NAND2X1 gate409 ( .A(N973), .B(N1470), .Y(N1501) );
  NAND2X1 gate410 ( .A(N994), .B(N1475), .Y(N1504) );
  INVX1 gate411 ( .A(N1464), .Y(N1510) );
  NAND2X1 gate412 ( .A(N1443), .B(N1487), .Y(N1513) );
  NAND2X1 gate413 ( .A(N1445), .B(N1488), .Y(N1514) );
  NAND2X1 gate414 ( .A(N1447), .B(N1489), .Y(N1517) );
  NAND2X1 gate415 ( .A(N1451), .B(N1492), .Y(N1520) );
  NAND2X1 gate416 ( .A(N1453), .B(N1493), .Y(N1521) );
  NAND2X1 gate417 ( .A(N1455), .B(N1494), .Y(N1522) );
  NAND2X1 gate418 ( .A(N1457), .B(N1495), .Y(N1526) );
  NAND2X1 gate419 ( .A(N1459), .B(N1496), .Y(N1527) );
  INVX1 gate420 ( .A(N1472), .Y(N1528) );
  NAND2X1 gate421 ( .A(N1462), .B(N1498), .Y(N1529) );
  INVX1 gate422 ( .A(N1478), .Y(N1530) );
  INVX1 gate423 ( .A(N1481), .Y(N1531) );
  INVX1 gate424 ( .A(N1484), .Y(N1532) );
  NAND2X1 gate425 ( .A(N1471), .B(N1501), .Y(N1534) );
  NAND2X1 gate426 ( .A(N1469), .B(N1500), .Y(N1537) );
  NAND2X1 gate427 ( .A(N1476), .B(N1504), .Y(N1540) );
  INVX1 gate428 ( .A(N1513), .Y(N1546) );
  INVX1 gate429 ( .A(N1521), .Y(N1554) );
  INVX1 gate430 ( .A(N1526), .Y(N1557) );
  INVX1 gate431 ( .A(N1520), .Y(N1561) );
  NAND2X1 gate432 ( .A(N1484), .B(N1531), .Y(N1567) );
  NAND2X1 gate433 ( .A(N1481), .B(N1532), .Y(N1568) );
  INVX1 gate434 ( .A(N1510), .Y(N1569) );
  INVX1 gate435 ( .A(N1527), .Y(N1571) );
  INVX1 gate436 ( .A(N1529), .Y(N1576) );
  BUFX2 gate437 ( .A(N1522), .Y(N1588) );
  INVX1 gate438 ( .A(N1534), .Y(N1591) );
  INVX1 gate439 ( .A(N1537), .Y(N1593) );
  NAND2X1 gate440 ( .A(N1540), .B(N1530), .Y(N1594) );
  INVX1 gate441 ( .A(N1540), .Y(N1595) );
  NAND2X1 gate442 ( .A(N1567), .B(N1568), .Y(N1596) );
  BUFX2 gate443 ( .A(N1517), .Y(N1600) );
  BUFX2 gate444 ( .A(N1517), .Y(N1603) );
  BUFX2 gate445 ( .A(N1522), .Y(N1606) );
  BUFX2 gate446 ( .A(N1522), .Y(N1609) );
  BUFX2 gate447 ( .A(N1514), .Y(N1612) );
  BUFX2 gate448 ( .A(N1514), .Y(N1615) );
  BUFX2 gate449 ( .A(N1557), .Y(N1620) );
  BUFX2 gate450 ( .A(N1554), .Y(N1623) );
  INVX1 gate451 ( .A(N1571), .Y(N1635) );
  NAND2X1 gate452 ( .A(N1478), .B(N1595), .Y(N1636) );
  NAND2X1 gate453 ( .A(N1576), .B(N1569), .Y(N1638) );
  INVX1 gate454 ( .A(N1576), .Y(N1639) );
  BUFX2 gate455 ( .A(N1561), .Y(N1640) );
  BUFX2 gate456 ( .A(N1561), .Y(N1643) );
  BUFX2 gate457 ( .A(N1546), .Y(N1647) );
  BUFX2 gate458 ( .A(N1546), .Y(N1651) );
  BUFX2 gate459 ( .A(N1554), .Y(N1658) );
  BUFX2 gate460 ( .A(N1557), .Y(N1661) );
  BUFX2 gate461 ( .A(N1557), .Y(N1664) );
  NAND2X1 gate462 ( .A(N1596), .B(N893), .Y(N1671) );
  INVX1 gate463 ( .A(N1596), .Y(N1672) );
  INVX1 gate464 ( .A(N1600), .Y(N1675) );
  INVX1 gate465 ( .A(N1603), .Y(N1677) );
  NAND2X1 gate466 ( .A(N1606), .B(N1217), .Y(N1678) );
  INVX1 gate467 ( .A(N1606), .Y(N1679) );
  NAND2X1 gate468 ( .A(N1609), .B(N1219), .Y(N1680) );
  INVX1 gate469 ( .A(N1609), .Y(N1681) );
  INVX1 gate470 ( .A(N1612), .Y(N1682) );
  INVX1 gate471 ( .A(N1615), .Y(N1683) );
  NAND2X1 gate472 ( .A(N1594), .B(N1636), .Y(N1685) );
  NAND2X1 gate473 ( .A(N1510), .B(N1639), .Y(N1688) );
  BUFX2 gate474 ( .A(N1588), .Y(N1697) );
  BUFX2 gate475 ( .A(N1588), .Y(N1701) );
  NAND2X1 gate476 ( .A(N643), .B(N1672), .Y(N1706) );
  INVX1 gate477 ( .A(N1643), .Y(N1707) );
  NAND2X1 gate478 ( .A(N1647), .B(N1675), .Y(N1708) );
  INVX1 gate479 ( .A(N1647), .Y(N1709) );
  NAND2X1 gate480 ( .A(N1651), .B(N1677), .Y(N1710) );
  INVX1 gate481 ( .A(N1651), .Y(N1711) );
  NAND2X1 gate482 ( .A(N1028), .B(N1679), .Y(N1712) );
  NAND2X1 gate483 ( .A(N1031), .B(N1681), .Y(N1713) );
  BUFX2 gate484 ( .A(N1620), .Y(N1714) );
  BUFX2 gate485 ( .A(N1620), .Y(N1717) );
  NAND2X1 gate486 ( .A(N1658), .B(N1593), .Y(N1720) );
  INVX1 gate487 ( .A(N1658), .Y(N1721) );
  NAND2X1 gate488 ( .A(N1638), .B(N1688), .Y(N1723) );
  INVX1 gate489 ( .A(N1661), .Y(N1727) );
  INVX1 gate490 ( .A(N1640), .Y(N1728) );
  INVX1 gate491 ( .A(N1664), .Y(N1730) );
  BUFX2 gate492 ( .A(N1623), .Y(N1731) );
  BUFX2 gate493 ( .A(N1623), .Y(N1734) );
  NAND2X1 gate494 ( .A(N1685), .B(N1528), .Y(N1740) );
  INVX1 gate495 ( .A(N1685), .Y(N1741) );
  NAND2X1 gate496 ( .A(N1671), .B(N1706), .Y(N1742) );
  NAND2X1 gate497 ( .A(N1600), .B(N1709), .Y(N1746) );
  NAND2X1 gate498 ( .A(N1603), .B(N1711), .Y(N1747) );
  NAND2X1 gate499 ( .A(N1678), .B(N1712), .Y(N1748) );
  NAND2X1 gate500 ( .A(N1680), .B(N1713), .Y(N1751) );
  NAND2X1 gate501 ( .A(N1537), .B(N1721), .Y(N1759) );
  INVX1 gate502 ( .A(N1697), .Y(N1761) );
  NAND2X1 gate503 ( .A(N1697), .B(N1727), .Y(N1762) );
  INVX1 gate504 ( .A(N1701), .Y(N1763) );
  NAND2X1 gate505 ( .A(N1701), .B(N1730), .Y(N1764) );
  INVX1 gate506 ( .A(N1717), .Y(N1768) );
  NAND2X1 gate507 ( .A(N1472), .B(N1741), .Y(N1769) );
  NAND2X1 gate508 ( .A(N1723), .B(N1413), .Y(N1772) );
  INVX1 gate509 ( .A(N1723), .Y(N1773) );
  NAND2X1 gate510 ( .A(N1708), .B(N1746), .Y(N1774) );
  NAND2X1 gate511 ( .A(N1710), .B(N1747), .Y(N1777) );
  INVX1 gate512 ( .A(N1731), .Y(N1783) );
  NAND2X1 gate513 ( .A(N1731), .B(N1682), .Y(N1784) );
  INVX1 gate514 ( .A(N1714), .Y(N1785) );
  INVX1 gate515 ( .A(N1734), .Y(N1786) );
  NAND2X1 gate516 ( .A(N1734), .B(N1683), .Y(N1787) );
  NAND2X1 gate517 ( .A(N1720), .B(N1759), .Y(N1788) );
  NAND2X1 gate518 ( .A(N1661), .B(N1761), .Y(N1791) );
  NAND2X1 gate519 ( .A(N1664), .B(N1763), .Y(N1792) );
  NAND2X1 gate520 ( .A(N1751), .B(N1155), .Y(N1795) );
  INVX1 gate521 ( .A(N1751), .Y(N1796) );
  NAND2X1 gate522 ( .A(N1740), .B(N1769), .Y(N1798) );
  NAND2X1 gate523 ( .A(N1334), .B(N1773), .Y(N1801) );
  NAND2X1 gate524 ( .A(N1742), .B(N290), .Y(N1802) );
  INVX1 gate525 ( .A(N1748), .Y(N1807) );
  NAND2X1 gate526 ( .A(N1748), .B(N1218), .Y(N1808) );
  NAND2X1 gate527 ( .A(N1612), .B(N1783), .Y(N1809) );
  NAND2X1 gate528 ( .A(N1615), .B(N1786), .Y(N1810) );
  NAND2X1 gate529 ( .A(N1791), .B(N1762), .Y(N1812) );
  NAND2X1 gate530 ( .A(N1792), .B(N1764), .Y(N1815) );
  BUFX2 gate531 ( .A(N1742), .Y(N1818) );
  NAND2X1 gate532 ( .A(N1777), .B(N1490), .Y(N1821) );
  INVX1 gate533 ( .A(N1777), .Y(N1822) );
  NAND2X1 gate534 ( .A(N1774), .B(N1491), .Y(N1823) );
  INVX1 gate535 ( .A(N1774), .Y(N1824) );
  NAND2X1 gate536 ( .A(N962), .B(N1796), .Y(N1825) );
  NAND2X1 gate537 ( .A(N1788), .B(N1409), .Y(N1826) );
  INVX1 gate538 ( .A(N1788), .Y(N1827) );
  NAND2X1 gate539 ( .A(N1772), .B(N1801), .Y(N1830) );
  NAND2X1 gate540 ( .A(N959), .B(N1807), .Y(N1837) );
  NAND2X1 gate541 ( .A(N1809), .B(N1784), .Y(N1838) );
  NAND2X1 gate542 ( .A(N1810), .B(N1787), .Y(N1841) );
  NAND2X1 gate543 ( .A(N1419), .B(N1822), .Y(N1848) );
  NAND2X1 gate544 ( .A(N1416), .B(N1824), .Y(N1849) );
  NAND2X1 gate545 ( .A(N1795), .B(N1825), .Y(N1850) );
  NAND2X1 gate546 ( .A(N1319), .B(N1827), .Y(N1852) );
  NAND2X1 gate547 ( .A(N1815), .B(N1707), .Y(N1855) );
  INVX1 gate548 ( .A(N1815), .Y(N1856) );
  INVX1 gate549 ( .A(N1818), .Y(N1857) );
  NAND2X1 gate550 ( .A(N1798), .B(N290), .Y(N1858) );
  INVX1 gate551 ( .A(N1812), .Y(N1864) );
  NAND2X1 gate552 ( .A(N1812), .B(N1728), .Y(N1865) );
  BUFX2 gate553 ( .A(N1798), .Y(N1866) );
  BUFX2 gate554 ( .A(N1802), .Y(N1869) );
  BUFX2 gate555 ( .A(N1802), .Y(N1872) );
  NAND2X1 gate556 ( .A(N1808), .B(N1837), .Y(N1875) );
  NAND2X1 gate557 ( .A(N1821), .B(N1848), .Y(N1878) );
  NAND2X1 gate558 ( .A(N1823), .B(N1849), .Y(N1879) );
  NAND2X1 gate559 ( .A(N1841), .B(N1768), .Y(N1882) );
  INVX1 gate560 ( .A(N1841), .Y(N1883) );
  NAND2X1 gate561 ( .A(N1826), .B(N1852), .Y(N1884) );
  NAND2X1 gate562 ( .A(N1643), .B(N1856), .Y(N1885) );
  NAND2X1 gate563 ( .A(N1830), .B(N290), .Y(N1889) );
  INVX1 gate564 ( .A(N1838), .Y(N1895) );
  NAND2X1 gate565 ( .A(N1838), .B(N1785), .Y(N1896) );
  NAND2X1 gate566 ( .A(N1640), .B(N1864), .Y(N1897) );
  INVX1 gate567 ( .A(N1850), .Y(N1898) );
  BUFX2 gate568 ( .A(N1830), .Y(N1902) );
  INVX1 gate569 ( .A(N1878), .Y(N1910) );
  NAND2X1 gate570 ( .A(N1717), .B(N1883), .Y(N1911) );
  INVX1 gate571 ( .A(N1884), .Y(N1912) );
  NAND2X1 gate572 ( .A(N1855), .B(N1885), .Y(N1913) );
  INVX1 gate573 ( .A(N1866), .Y(N1915) );
  NAND2X1 gate574 ( .A(N1872), .B(N919), .Y(N1919) );
  INVX1 gate575 ( .A(N1872), .Y(N1920) );
  NAND2X1 gate576 ( .A(N1869), .B(N920), .Y(N1921) );
  INVX1 gate577 ( .A(N1869), .Y(N1922) );
  INVX1 gate578 ( .A(N1875), .Y(N1923) );
  NAND2X1 gate579 ( .A(N1714), .B(N1895), .Y(N1924) );
  BUFX2 gate580 ( .A(N1858), .Y(N1927) );
  BUFX2 gate581 ( .A(N1858), .Y(N1930) );
  NAND2X1 gate582 ( .A(N1865), .B(N1897), .Y(N1933) );
  NAND2X1 gate583 ( .A(N1882), .B(N1911), .Y(N1936) );
  INVX1 gate584 ( .A(N1898), .Y(N1937) );
  INVX1 gate585 ( .A(N1902), .Y(N1938) );
  NAND2X1 gate586 ( .A(N679), .B(N1920), .Y(N1941) );
  NAND2X1 gate587 ( .A(N676), .B(N1922), .Y(N1942) );
  BUFX2 gate588 ( .A(N1879), .Y(N1944) );
  INVX1 gate589 ( .A(N1913), .Y(N1947) );
  BUFX2 gate590 ( .A(N1889), .Y(N1950) );
  BUFX2 gate591 ( .A(N1889), .Y(N1953) );
  BUFX2 gate592 ( .A(N1879), .Y(N1958) );
  NAND2X1 gate593 ( .A(N1896), .B(N1924), .Y(N1961) );
  AND2X1 gate594 ( .A(N1910), .B(N601), .Y(N1965) );
  AND2X1 gate595 ( .A(N602), .B(N1912), .Y(N1968) );
  NAND2X1 gate596 ( .A(N1930), .B(N917), .Y(N1975) );
  INVX1 gate597 ( .A(N1930), .Y(N1976) );
  NAND2X1 gate598 ( .A(N1927), .B(N918), .Y(N1977) );
  INVX1 gate599 ( .A(N1927), .Y(N1978) );
  NAND2X1 gate600 ( .A(N1919), .B(N1941), .Y(N1979) );
  NAND2X1 gate601 ( .A(N1921), .B(N1942), .Y(N1980) );
  INVX1 gate602 ( .A(N1933), .Y(N1985) );
  INVX1 gate603 ( .A(N1936), .Y(N1987) );
  INVX1 gate604 ( .A(N1944), .Y(N1999) );
  NAND2X1 gate605 ( .A(N1944), .B(N1937), .Y(N2000) );
  INVX1 gate606 ( .A(N1947), .Y(N2002) );
  NAND2X1 gate607 ( .A(N1947), .B(N1499), .Y(N2003) );
  NAND2X1 gate608 ( .A(N1953), .B(N1350), .Y(N2004) );
  INVX1 gate609 ( .A(N1953), .Y(N2005) );
  NAND2X1 gate610 ( .A(N1950), .B(N1351), .Y(N2006) );
  INVX1 gate611 ( .A(N1950), .Y(N2007) );
  NAND2X1 gate612 ( .A(N673), .B(N1976), .Y(N2008) );
  NAND2X1 gate613 ( .A(N670), .B(N1978), .Y(N2009) );
  INVX1 gate614 ( .A(N1979), .Y(N2012) );
  INVX1 gate615 ( .A(N1958), .Y(N2013) );
  NAND2X1 gate616 ( .A(N1958), .B(N1923), .Y(N2014) );
  INVX1 gate617 ( .A(N1961), .Y(N2015) );
  NAND2X1 gate618 ( .A(N1961), .B(N1635), .Y(N2016) );
  INVX1 gate619 ( .A(N1965), .Y(N2018) );
  INVX1 gate620 ( .A(N1968), .Y(N2019) );
  NAND2X1 gate621 ( .A(N1898), .B(N1999), .Y(N2020) );
  INVX1 gate622 ( .A(N1987), .Y(N2021) );
  NAND2X1 gate623 ( .A(N1987), .B(N1591), .Y(N2022) );
  NAND2X1 gate624 ( .A(N1440), .B(N2002), .Y(N2023) );
  NAND2X1 gate625 ( .A(N1261), .B(N2005), .Y(N2024) );
  NAND2X1 gate626 ( .A(N1258), .B(N2007), .Y(N2025) );
  NAND2X1 gate627 ( .A(N1975), .B(N2008), .Y(N2026) );
  NAND2X1 gate628 ( .A(N1977), .B(N2009), .Y(N2027) );
  INVX1 gate629 ( .A(N1980), .Y(N2030) );
  BUFX2 gate630 ( .A(N1980), .Y(N2033) );
  NAND2X1 gate631 ( .A(N1875), .B(N2013), .Y(N2036) );
  NAND2X1 gate632 ( .A(N1571), .B(N2015), .Y(N2037) );
  NAND2X1 gate633 ( .A(N2020), .B(N2000), .Y(N2038) );
  NAND2X1 gate634 ( .A(N1534), .B(N2021), .Y(N2039) );
  NAND2X1 gate635 ( .A(N2023), .B(N2003), .Y(N2040) );
  NAND2X1 gate636 ( .A(N2004), .B(N2024), .Y(N2041) );
  NAND2X1 gate637 ( .A(N2006), .B(N2025), .Y(N2042) );
  INVX1 gate638 ( .A(N2026), .Y(N2047) );
  NAND2X1 gate639 ( .A(N2036), .B(N2014), .Y(N2052) );
  NAND2X1 gate640 ( .A(N2037), .B(N2016), .Y(N2055) );
  INVX1 gate641 ( .A(N2038), .Y(N2060) );
  NAND2X1 gate642 ( .A(N2039), .B(N2022), .Y(N2061) );
  NAND2X1 gate643 ( .A(N2040), .B(N290), .Y(N2062) );
  INVX1 gate644 ( .A(N2041), .Y(N2067) );
  INVX1 gate645 ( .A(N2027), .Y(N2068) );
  BUFX2 gate646 ( .A(N2027), .Y(N2071) );
  INVX1 gate647 ( .A(N2052), .Y(N2076) );
  INVX1 gate648 ( .A(N2055), .Y(N2077) );
  NAND2X1 gate649 ( .A(N2060), .B(N290), .Y(N2078) );
  NAND2X1 gate650 ( .A(N2061), .B(N290), .Y(N2081) );
  INVX1 gate651 ( .A(N2042), .Y(N2086) );
  BUFX2 gate652 ( .A(N2042), .Y(N2089) );
  AND2X1 gate653 ( .A(N2030), .B(N2068), .Y(N2104) );
  AND2X1 gate654 ( .A(N2033), .B(N2068), .Y(N2119) );
  AND2X1 gate655 ( .A(N2030), .B(N2071), .Y(N2129) );
  AND2X1 gate656 ( .A(N2033), .B(N2071), .Y(N2143) );
  BUFX2 gate657 ( .A(N2062), .Y(N2148) );
  BUFX2 gate658 ( .A(N2062), .Y(N2151) );
  BUFX2 gate659 ( .A(N2078), .Y(N2196) );
  BUFX2 gate660 ( .A(N2078), .Y(N2199) );
  BUFX2 gate661 ( .A(N2081), .Y(N2202) );
  BUFX2 gate662 ( .A(N2081), .Y(N2205) );
  NAND2X1 gate663 ( .A(N2151), .B(N915), .Y(N2214) );
  INVX1 gate664 ( .A(N2151), .Y(N2215) );
  NAND2X1 gate665 ( .A(N2148), .B(N916), .Y(N2216) );
  INVX1 gate666 ( .A(N2148), .Y(N2217) );
  NAND2X1 gate667 ( .A(N2199), .B(N1348), .Y(N2222) );
  INVX1 gate668 ( .A(N2199), .Y(N2223) );
  NAND2X1 gate669 ( .A(N2196), .B(N1349), .Y(N2224) );
  INVX1 gate670 ( .A(N2196), .Y(N2225) );
  NAND2X1 gate671 ( .A(N2205), .B(N913), .Y(N2226) );
  INVX1 gate672 ( .A(N2205), .Y(N2227) );
  NAND2X1 gate673 ( .A(N2202), .B(N914), .Y(N2228) );
  INVX1 gate674 ( .A(N2202), .Y(N2229) );
  NAND2X1 gate675 ( .A(N667), .B(N2215), .Y(N2230) );
  NAND2X1 gate676 ( .A(N664), .B(N2217), .Y(N2231) );
  NAND2X1 gate677 ( .A(N1255), .B(N2223), .Y(N2232) );
  NAND2X1 gate678 ( .A(N1252), .B(N2225), .Y(N2233) );
  NAND2X1 gate679 ( .A(N661), .B(N2227), .Y(N2234) );
  NAND2X1 gate680 ( .A(N658), .B(N2229), .Y(N2235) );
  NAND2X1 gate681 ( .A(N2214), .B(N2230), .Y(N2236) );
  NAND2X1 gate682 ( .A(N2216), .B(N2231), .Y(N2237) );
  NAND2X1 gate683 ( .A(N2222), .B(N2232), .Y(N2240) );
  NAND2X1 gate684 ( .A(N2224), .B(N2233), .Y(N2241) );
  NAND2X1 gate685 ( .A(N2226), .B(N2234), .Y(N2244) );
  NAND2X1 gate686 ( .A(N2228), .B(N2235), .Y(N2245) );
  INVX1 gate687 ( .A(N2236), .Y(N2250) );
  INVX1 gate688 ( .A(N2240), .Y(N2253) );
  INVX1 gate689 ( .A(N2244), .Y(N2256) );
  INVX1 gate690 ( .A(N2237), .Y(N2257) );
  BUFX2 gate691 ( .A(N2237), .Y(N2260) );
  INVX1 gate692 ( .A(N2241), .Y(N2263) );
  AND2X1 gate693 ( .A(N1164), .B(N2241), .Y(N2266) );
  INVX1 gate694 ( .A(N2245), .Y(N2269) );
  AND2X1 gate695 ( .A(N1168), .B(N2245), .Y(N2272) );
  NAND3X1 gate696_1 ( .A(N2067), .B(N2012), .C(N2047), .Y(N2279_1) );
  NAND3X1 gate696_2 ( .A(N2250), .B(N899), .C(N2256), .Y(N2279_2) );
  NAND3X1 gate696_3 ( .A(N2253), .B(N903), .C(N2279_1), .Y(N2279_3) );
  NAND2X1 gate696 ( .A(N2279_2), .B(N2279_3), .Y(N2279) );
  BUFX2 gate697 ( .A(N2266), .Y(N2286) );
  BUFX2 gate698 ( .A(N2266), .Y(N2297) );
  BUFX2 gate699 ( .A(N2272), .Y(N2315) );
  BUFX2 gate700 ( .A(N2272), .Y(N2326) );
  AND2X1 gate701 ( .A(N2086), .B(N2257), .Y(N2340) );
  AND2X1 gate702 ( .A(N2089), .B(N2257), .Y(N2353) );
  AND2X1 gate703 ( .A(N2086), .B(N2260), .Y(N2361) );
  AND2X1 gate704 ( .A(N2089), .B(N2260), .Y(N2375) );
  AND2X1 gate705_1 ( .A(N338), .B(N2279), .Y(N2384_1) );
  AND2X1 gate705_2 ( .A(N313), .B(N313), .Y(N2384_2) );
  AND2X1 gate705 ( .A(N2384_1), .B(N2384_2), .Y(N2384) );
  AND2X1 gate706 ( .A(N1163), .B(N2263), .Y(N2385) );
  AND2X1 gate707 ( .A(N1164), .B(N2263), .Y(N2386) );
  AND2X1 gate708 ( .A(N1167), .B(N2269), .Y(N2426) );
  AND2X1 gate709 ( .A(N1168), .B(N2269), .Y(N2427) );
  NAND3X1 gate710_1 ( .A(N2286), .B(N2315), .C(N2361), .Y(N2537_1) );
  NAND2X1 gate710_2 ( .A(N2104), .B(N1171), .Y(N2537_2) );
  NAND2X1 gate710 ( .A(N2537_1), .B(N2537_2), .Y(N2537) );
  NAND3X1 gate711_1 ( .A(N2286), .B(N2315), .C(N2340), .Y(N2540_1) );
  NAND2X1 gate711_2 ( .A(N2129), .B(N1171), .Y(N2540_2) );
  NAND2X1 gate711 ( .A(N2540_1), .B(N2540_2), .Y(N2540) );
  NAND3X1 gate712_1 ( .A(N2286), .B(N2315), .C(N2340), .Y(N2543_1) );
  NAND2X1 gate712_2 ( .A(N2119), .B(N1171), .Y(N2543_2) );
  NAND2X1 gate712 ( .A(N2543_1), .B(N2543_2), .Y(N2543) );
  NAND3X1 gate713_1 ( .A(N2286), .B(N2315), .C(N2353), .Y(N2546_1) );
  NAND2X1 gate713_2 ( .A(N2104), .B(N1171), .Y(N2546_2) );
  NAND2X1 gate713 ( .A(N2546_1), .B(N2546_2), .Y(N2546) );
  NAND3X1 gate714_1 ( .A(N2297), .B(N2315), .C(N2375), .Y(N2549_1) );
  NAND2X1 gate714_2 ( .A(N2119), .B(N1188), .Y(N2549_2) );
  NAND2X1 gate714 ( .A(N2549_1), .B(N2549_2), .Y(N2549) );
  NAND3X1 gate715_1 ( .A(N2297), .B(N2326), .C(N2361), .Y(N2552_1) );
  NAND2X1 gate715_2 ( .A(N2143), .B(N1188), .Y(N2552_2) );
  NAND2X1 gate715 ( .A(N2552_1), .B(N2552_2), .Y(N2552) );
  NAND3X1 gate716_1 ( .A(N2297), .B(N2326), .C(N2375), .Y(N2555_1) );
  NAND2X1 gate716_2 ( .A(N2129), .B(N1188), .Y(N2555_2) );
  NAND2X1 gate716 ( .A(N2555_1), .B(N2555_2), .Y(N2555) );
  AND2X1 gate717_1 ( .A(N2286), .B(N2315), .Y(N2558_1) );
  AND2X1 gate717_2 ( .A(N2361), .B(N2104), .Y(N2558_2) );
  AND2X1 gate717_3 ( .A(N1171), .B(N2558_1), .Y(N2558_3) );
  AND2X1 gate717 ( .A(N2558_2), .B(N2558_3), .Y(N2558) );
  AND2X1 gate718_1 ( .A(N2286), .B(N2315), .Y(N2561_1) );
  AND2X1 gate718_2 ( .A(N2340), .B(N2129), .Y(N2561_2) );
  AND2X1 gate718_3 ( .A(N1171), .B(N2561_1), .Y(N2561_3) );
  AND2X1 gate718 ( .A(N2561_2), .B(N2561_3), .Y(N2561) );
  AND2X1 gate719_1 ( .A(N2286), .B(N2315), .Y(N2564_1) );
  AND2X1 gate719_2 ( .A(N2340), .B(N2119), .Y(N2564_2) );
  AND2X1 gate719_3 ( .A(N1171), .B(N2564_1), .Y(N2564_3) );
  AND2X1 gate719 ( .A(N2564_2), .B(N2564_3), .Y(N2564) );
  AND2X1 gate720_1 ( .A(N2286), .B(N2315), .Y(N2567_1) );
  AND2X1 gate720_2 ( .A(N2353), .B(N2104), .Y(N2567_2) );
  AND2X1 gate720_3 ( .A(N1171), .B(N2567_1), .Y(N2567_3) );
  AND2X1 gate720 ( .A(N2567_2), .B(N2567_3), .Y(N2567) );
  AND2X1 gate721_1 ( .A(N2297), .B(N2315), .Y(N2570_1) );
  AND2X1 gate721_2 ( .A(N2375), .B(N2119), .Y(N2570_2) );
  AND2X1 gate721_3 ( .A(N1188), .B(N2570_1), .Y(N2570_3) );
  AND2X1 gate721 ( .A(N2570_2), .B(N2570_3), .Y(N2570) );
  AND2X1 gate722_1 ( .A(N2297), .B(N2326), .Y(N2573_1) );
  AND2X1 gate722_2 ( .A(N2361), .B(N2143), .Y(N2573_2) );
  AND2X1 gate722_3 ( .A(N1188), .B(N2573_1), .Y(N2573_3) );
  AND2X1 gate722 ( .A(N2573_2), .B(N2573_3), .Y(N2573) );
  AND2X1 gate723_1 ( .A(N2297), .B(N2326), .Y(N2576_1) );
  AND2X1 gate723_2 ( .A(N2375), .B(N2129), .Y(N2576_2) );
  AND2X1 gate723_3 ( .A(N1188), .B(N2576_1), .Y(N2576_3) );
  AND2X1 gate723 ( .A(N2576_2), .B(N2576_3), .Y(N2576) );
  NAND3X1 gate724_1 ( .A(N2286), .B(N2427), .C(N2361), .Y(N2594_1) );
  NAND2X1 gate724_2 ( .A(N2129), .B(N1171), .Y(N2594_2) );
  NAND2X1 gate724 ( .A(N2594_1), .B(N2594_2), .Y(N2594) );
  NAND3X1 gate725_1 ( .A(N2297), .B(N2427), .C(N2361), .Y(N2597_1) );
  NAND2X1 gate725_2 ( .A(N2119), .B(N1171), .Y(N2597_2) );
  NAND2X1 gate725 ( .A(N2597_1), .B(N2597_2), .Y(N2597) );
  NAND3X1 gate726_1 ( .A(N2297), .B(N2427), .C(N2375), .Y(N2600_1) );
  NAND2X1 gate726_2 ( .A(N2104), .B(N1171), .Y(N2600_2) );
  NAND2X1 gate726 ( .A(N2600_1), .B(N2600_2), .Y(N2600) );
  NAND3X1 gate727_1 ( .A(N2297), .B(N2427), .C(N2340), .Y(N2603_1) );
  NAND2X1 gate727_2 ( .A(N2143), .B(N1171), .Y(N2603_2) );
  NAND2X1 gate727 ( .A(N2603_1), .B(N2603_2), .Y(N2603) );
  NAND3X1 gate728_1 ( .A(N2297), .B(N2427), .C(N2353), .Y(N2606_1) );
  NAND2X1 gate728_2 ( .A(N2129), .B(N1188), .Y(N2606_2) );
  NAND2X1 gate728 ( .A(N2606_1), .B(N2606_2), .Y(N2606) );
  NAND3X1 gate729_1 ( .A(N2386), .B(N2326), .C(N2361), .Y(N2611_1) );
  NAND2X1 gate729_2 ( .A(N2129), .B(N1188), .Y(N2611_2) );
  NAND2X1 gate729 ( .A(N2611_1), .B(N2611_2), .Y(N2611) );
  NAND3X1 gate730_1 ( .A(N2386), .B(N2326), .C(N2361), .Y(N2614_1) );
  NAND2X1 gate730_2 ( .A(N2119), .B(N1188), .Y(N2614_2) );
  NAND2X1 gate730 ( .A(N2614_1), .B(N2614_2), .Y(N2614) );
  NAND3X1 gate731_1 ( .A(N2386), .B(N2326), .C(N2375), .Y(N2617_1) );
  NAND2X1 gate731_2 ( .A(N2104), .B(N1188), .Y(N2617_2) );
  NAND2X1 gate731 ( .A(N2617_1), .B(N2617_2), .Y(N2617) );
  NAND3X1 gate732_1 ( .A(N2386), .B(N2326), .C(N2353), .Y(N2620_1) );
  NAND2X1 gate732_2 ( .A(N2129), .B(N1188), .Y(N2620_2) );
  NAND2X1 gate732 ( .A(N2620_1), .B(N2620_2), .Y(N2620) );
  NAND3X1 gate733_1 ( .A(N2297), .B(N2427), .C(N2340), .Y(N2627_1) );
  NAND2X1 gate733_2 ( .A(N2104), .B(N926), .Y(N2627_2) );
  NAND2X1 gate733 ( .A(N2627_1), .B(N2627_2), .Y(N2627) );
  NAND3X1 gate734_1 ( .A(N2386), .B(N2326), .C(N2340), .Y(N2628_1) );
  NAND2X1 gate734_2 ( .A(N2104), .B(N926), .Y(N2628_2) );
  NAND2X1 gate734 ( .A(N2628_1), .B(N2628_2), .Y(N2628) );
  NAND3X1 gate735_1 ( .A(N2386), .B(N2427), .C(N2361), .Y(N2629_1) );
  NAND2X1 gate735_2 ( .A(N2104), .B(N926), .Y(N2629_2) );
  NAND2X1 gate735 ( .A(N2629_1), .B(N2629_2), .Y(N2629) );
  NAND3X1 gate736_1 ( .A(N2386), .B(N2427), .C(N2340), .Y(N2630_1) );
  NAND2X1 gate736_2 ( .A(N2129), .B(N926), .Y(N2630_2) );
  NAND2X1 gate736 ( .A(N2630_1), .B(N2630_2), .Y(N2630) );
  NAND3X1 gate737_1 ( .A(N2386), .B(N2427), .C(N2340), .Y(N2631_1) );
  NAND2X1 gate737_2 ( .A(N2119), .B(N926), .Y(N2631_2) );
  NAND2X1 gate737 ( .A(N2631_1), .B(N2631_2), .Y(N2631) );
  NAND3X1 gate738_1 ( .A(N2386), .B(N2427), .C(N2353), .Y(N2632_1) );
  NAND2X1 gate738_2 ( .A(N2104), .B(N926), .Y(N2632_2) );
  NAND2X1 gate738 ( .A(N2632_1), .B(N2632_2), .Y(N2632) );
  NAND3X1 gate739_1 ( .A(N2386), .B(N2426), .C(N2340), .Y(N2633_1) );
  NAND2X1 gate739_2 ( .A(N2104), .B(N926), .Y(N2633_2) );
  NAND2X1 gate739 ( .A(N2633_1), .B(N2633_2), .Y(N2633) );
  NAND3X1 gate740_1 ( .A(N2385), .B(N2427), .C(N2340), .Y(N2634_1) );
  NAND2X1 gate740_2 ( .A(N2104), .B(N926), .Y(N2634_2) );
  NAND2X1 gate740 ( .A(N2634_1), .B(N2634_2), .Y(N2634) );
  AND2X1 gate741_1 ( .A(N2286), .B(N2427), .Y(N2639_1) );
  AND2X1 gate741_2 ( .A(N2361), .B(N2129), .Y(N2639_2) );
  AND2X1 gate741_3 ( .A(N1171), .B(N2639_1), .Y(N2639_3) );
  AND2X1 gate741 ( .A(N2639_2), .B(N2639_3), .Y(N2639) );
  AND2X1 gate742_1 ( .A(N2297), .B(N2427), .Y(N2642_1) );
  AND2X1 gate742_2 ( .A(N2361), .B(N2119), .Y(N2642_2) );
  AND2X1 gate742_3 ( .A(N1171), .B(N2642_1), .Y(N2642_3) );
  AND2X1 gate742 ( .A(N2642_2), .B(N2642_3), .Y(N2642) );
  AND2X1 gate743_1 ( .A(N2297), .B(N2427), .Y(N2645_1) );
  AND2X1 gate743_2 ( .A(N2375), .B(N2104), .Y(N2645_2) );
  AND2X1 gate743_3 ( .A(N1171), .B(N2645_1), .Y(N2645_3) );
  AND2X1 gate743 ( .A(N2645_2), .B(N2645_3), .Y(N2645) );
  AND2X1 gate744_1 ( .A(N2297), .B(N2427), .Y(N2648_1) );
  AND2X1 gate744_2 ( .A(N2340), .B(N2143), .Y(N2648_2) );
  AND2X1 gate744_3 ( .A(N1171), .B(N2648_1), .Y(N2648_3) );
  AND2X1 gate744 ( .A(N2648_2), .B(N2648_3), .Y(N2648) );
  AND2X1 gate745_1 ( .A(N2297), .B(N2427), .Y(N2651_1) );
  AND2X1 gate745_2 ( .A(N2353), .B(N2129), .Y(N2651_2) );
  AND2X1 gate745_3 ( .A(N1188), .B(N2651_1), .Y(N2651_3) );
  AND2X1 gate745 ( .A(N2651_2), .B(N2651_3), .Y(N2651) );
  AND2X1 gate746_1 ( .A(N2386), .B(N2326), .Y(N2655_1) );
  AND2X1 gate746_2 ( .A(N2361), .B(N2129), .Y(N2655_2) );
  AND2X1 gate746_3 ( .A(N1188), .B(N2655_1), .Y(N2655_3) );
  AND2X1 gate746 ( .A(N2655_2), .B(N2655_3), .Y(N2655) );
  AND2X1 gate747_1 ( .A(N2386), .B(N2326), .Y(N2658_1) );
  AND2X1 gate747_2 ( .A(N2361), .B(N2119), .Y(N2658_2) );
  AND2X1 gate747_3 ( .A(N1188), .B(N2658_1), .Y(N2658_3) );
  AND2X1 gate747 ( .A(N2658_2), .B(N2658_3), .Y(N2658) );
  AND2X1 gate748_1 ( .A(N2386), .B(N2326), .Y(N2661_1) );
  AND2X1 gate748_2 ( .A(N2375), .B(N2104), .Y(N2661_2) );
  AND2X1 gate748_3 ( .A(N1188), .B(N2661_1), .Y(N2661_3) );
  AND2X1 gate748 ( .A(N2661_2), .B(N2661_3), .Y(N2661) );
  AND2X1 gate749_1 ( .A(N2386), .B(N2326), .Y(N2664_1) );
  AND2X1 gate749_2 ( .A(N2353), .B(N2129), .Y(N2664_2) );
  AND2X1 gate749_3 ( .A(N1188), .B(N2664_1), .Y(N2664_3) );
  AND2X1 gate749 ( .A(N2664_2), .B(N2664_3), .Y(N2664) );
  NAND2X1 gate750 ( .A(N2558), .B(N534), .Y(N2669) );
  INVX1 gate751 ( .A(N2558), .Y(N2670) );
  NAND2X1 gate752 ( .A(N2561), .B(N535), .Y(N2671) );
  INVX1 gate753 ( .A(N2561), .Y(N2672) );
  NAND2X1 gate754 ( .A(N2564), .B(N536), .Y(N2673) );
  INVX1 gate755 ( .A(N2564), .Y(N2674) );
  NAND2X1 gate756 ( .A(N2567), .B(N537), .Y(N2675) );
  INVX1 gate757 ( .A(N2567), .Y(N2676) );
  NAND2X1 gate758 ( .A(N2570), .B(N543), .Y(N2682) );
  INVX1 gate759 ( .A(N2570), .Y(N2683) );
  NAND2X1 gate760 ( .A(N2573), .B(N548), .Y(N2688) );
  INVX1 gate761 ( .A(N2573), .Y(N2689) );
  NAND2X1 gate762 ( .A(N2576), .B(N549), .Y(N2690) );
  INVX1 gate763 ( .A(N2576), .Y(N2691) );
  AND2X1 gate764_1 ( .A(N2627), .B(N2628), .Y(N2710_1) );
  AND2X1 gate764_2 ( .A(N2629), .B(N2630), .Y(N2710_2) );
  AND2X1 gate764_3 ( .A(N2631), .B(N2632), .Y(N2710_3) );
  AND2X1 gate764_4 ( .A(N2633), .B(N2634), .Y(N2710_4) );
  AND2X1 gate764_5 ( .A(N2710_1), .B(N2710_2), .Y(N2710_5) );
  AND2X1 gate764_6 ( .A(N2710_3), .B(N2710_4), .Y(N2710_6) );
  AND2X1 gate764 ( .A(N2710_5), .B(N2710_6), .Y(N2710) );
  NAND2X1 gate765 ( .A(N343), .B(N2670), .Y(N2720) );
  NAND2X1 gate766 ( .A(N346), .B(N2672), .Y(N2721) );
  NAND2X1 gate767 ( .A(N349), .B(N2674), .Y(N2722) );
  NAND2X1 gate768 ( .A(N352), .B(N2676), .Y(N2723) );
  NAND2X1 gate769 ( .A(N2639), .B(N538), .Y(N2724) );
  INVX1 gate770 ( .A(N2639), .Y(N2725) );
  NAND2X1 gate771 ( .A(N2642), .B(N539), .Y(N2726) );
  INVX1 gate772 ( .A(N2642), .Y(N2727) );
  NAND2X1 gate773 ( .A(N2645), .B(N540), .Y(N2728) );
  INVX1 gate774 ( .A(N2645), .Y(N2729) );
  NAND2X1 gate775 ( .A(N2648), .B(N541), .Y(N2730) );
  INVX1 gate776 ( .A(N2648), .Y(N2731) );
  NAND2X1 gate777 ( .A(N2651), .B(N542), .Y(N2732) );
  INVX1 gate778 ( .A(N2651), .Y(N2733) );
  NAND2X1 gate779 ( .A(N370), .B(N2683), .Y(N2734) );
  NAND2X1 gate780 ( .A(N2655), .B(N544), .Y(N2735) );
  INVX1 gate781 ( .A(N2655), .Y(N2736) );
  NAND2X1 gate782 ( .A(N2658), .B(N545), .Y(N2737) );
  INVX1 gate783 ( .A(N2658), .Y(N2738) );
  NAND2X1 gate784 ( .A(N2661), .B(N546), .Y(N2739) );
  INVX1 gate785 ( .A(N2661), .Y(N2740) );
  NAND2X1 gate786 ( .A(N2664), .B(N547), .Y(N2741) );
  INVX1 gate787 ( .A(N2664), .Y(N2742) );
  NAND2X1 gate788 ( .A(N385), .B(N2689), .Y(N2743) );
  NAND2X1 gate789 ( .A(N388), .B(N2691), .Y(N2744) );
  NAND3X1 gate790_1 ( .A(N2537), .B(N2540), .C(N2543), .Y(N2745_1) );
  NAND3X1 gate790_2 ( .A(N2546), .B(N2594), .C(N2597), .Y(N2745_2) );
  NAND3X1 gate790_3 ( .A(N2600), .B(N2603), .C(N2745_1), .Y(N2745_3) );
  NAND2X1 gate790 ( .A(N2745_2), .B(N2745_3), .Y(N2745) );
  NAND3X1 gate791_1 ( .A(N2606), .B(N2549), .C(N2611), .Y(N2746_1) );
  NAND3X1 gate791_2 ( .A(N2614), .B(N2617), .C(N2620), .Y(N2746_2) );
  NAND3X1 gate791_3 ( .A(N2552), .B(N2555), .C(N2746_1), .Y(N2746_3) );
  NAND2X1 gate791 ( .A(N2746_2), .B(N2746_3), .Y(N2746) );
  AND2X1 gate792_1 ( .A(N2537), .B(N2540), .Y(N2747_1) );
  AND2X1 gate792_2 ( .A(N2543), .B(N2546), .Y(N2747_2) );
  AND2X1 gate792_3 ( .A(N2594), .B(N2597), .Y(N2747_3) );
  AND2X1 gate792_4 ( .A(N2600), .B(N2603), .Y(N2747_4) );
  AND2X1 gate792_5 ( .A(N2747_1), .B(N2747_2), .Y(N2747_5) );
  AND2X1 gate792_6 ( .A(N2747_3), .B(N2747_4), .Y(N2747_6) );
  AND2X1 gate792 ( .A(N2747_5), .B(N2747_6), .Y(N2747) );
  AND2X1 gate793_1 ( .A(N2606), .B(N2549), .Y(N2750_1) );
  AND2X1 gate793_2 ( .A(N2611), .B(N2614), .Y(N2750_2) );
  AND2X1 gate793_3 ( .A(N2617), .B(N2620), .Y(N2750_3) );
  AND2X1 gate793_4 ( .A(N2552), .B(N2555), .Y(N2750_4) );
  AND2X1 gate793_5 ( .A(N2750_1), .B(N2750_2), .Y(N2750_5) );
  AND2X1 gate793_6 ( .A(N2750_3), .B(N2750_4), .Y(N2750_6) );
  AND2X1 gate793 ( .A(N2750_5), .B(N2750_6), .Y(N2750) );
  NAND2X1 gate794 ( .A(N2669), .B(N2720), .Y(N2753) );
  NAND2X1 gate795 ( .A(N2671), .B(N2721), .Y(N2754) );
  NAND2X1 gate796 ( .A(N2673), .B(N2722), .Y(N2755) );
  NAND2X1 gate797 ( .A(N2675), .B(N2723), .Y(N2756) );
  NAND2X1 gate798 ( .A(N355), .B(N2725), .Y(N2757) );
  NAND2X1 gate799 ( .A(N358), .B(N2727), .Y(N2758) );
  NAND2X1 gate800 ( .A(N361), .B(N2729), .Y(N2759) );
  NAND2X1 gate801 ( .A(N364), .B(N2731), .Y(N2760) );
  NAND2X1 gate802 ( .A(N367), .B(N2733), .Y(N2761) );
  NAND2X1 gate803 ( .A(N2682), .B(N2734), .Y(N2762) );
  NAND2X1 gate804 ( .A(N373), .B(N2736), .Y(N2763) );
  NAND2X1 gate805 ( .A(N376), .B(N2738), .Y(N2764) );
  NAND2X1 gate806 ( .A(N379), .B(N2740), .Y(N2765) );
  NAND2X1 gate807 ( .A(N382), .B(N2742), .Y(N2766) );
  NAND2X1 gate808 ( .A(N2688), .B(N2743), .Y(N2767) );
  NAND2X1 gate809 ( .A(N2690), .B(N2744), .Y(N2768) );
  AND2X1 gate810 ( .A(N2745), .B(N275), .Y(N2773) );
  AND2X1 gate811 ( .A(N2746), .B(N276), .Y(N2776) );
  NAND2X1 gate812 ( .A(N2724), .B(N2757), .Y(N2779) );
  NAND2X1 gate813 ( .A(N2726), .B(N2758), .Y(N2780) );
  NAND2X1 gate814 ( .A(N2728), .B(N2759), .Y(N2781) );
  NAND2X1 gate815 ( .A(N2730), .B(N2760), .Y(N2782) );
  NAND2X1 gate816 ( .A(N2732), .B(N2761), .Y(N2783) );
  NAND2X1 gate817 ( .A(N2735), .B(N2763), .Y(N2784) );
  NAND2X1 gate818 ( .A(N2737), .B(N2764), .Y(N2785) );
  NAND2X1 gate819 ( .A(N2739), .B(N2765), .Y(N2786) );
  NAND2X1 gate820 ( .A(N2741), .B(N2766), .Y(N2787) );
  AND2X1 gate821_1 ( .A(N2747), .B(N2750), .Y(N2788_1) );
  AND2X1 gate821 ( .A(N2710), .B(N2788_1), .Y(N2788) );
  NAND2X1 gate822 ( .A(N2747), .B(N2750), .Y(N2789) );
  AND2X1 gate823_1 ( .A(N338), .B(N2279), .Y(N2800_1) );
  AND2X1 gate823_2 ( .A(N99), .B(N2788), .Y(N2800_2) );
  AND2X1 gate823 ( .A(N2800_1), .B(N2800_2), .Y(N2800) );
  NAND2X1 gate824 ( .A(N2773), .B(N2018), .Y(N2807) );
  INVX1 gate825 ( .A(N2773), .Y(N2808) );
  NAND2X1 gate826 ( .A(N2776), .B(N2019), .Y(N2809) );
  INVX1 gate827 ( .A(N2776), .Y(N2810) );
  NOR2X1 gate828 ( .A(N2384), .B(N2800), .Y(N2811) );
  AND2X1 gate829_1 ( .A(N897), .B(N283), .Y(N2812_1) );
  AND2X1 gate829 ( .A(N2789), .B(N2812_1), .Y(N2812) );
  AND2X1 gate830_1 ( .A(N76), .B(N283), .Y(N2815_1) );
  AND2X1 gate830 ( .A(N2789), .B(N2815_1), .Y(N2815) );
  AND2X1 gate831_1 ( .A(N82), .B(N283), .Y(N2818_1) );
  AND2X1 gate831 ( .A(N2789), .B(N2818_1), .Y(N2818) );
  AND2X1 gate832_1 ( .A(N85), .B(N283), .Y(N2821_1) );
  AND2X1 gate832 ( .A(N2789), .B(N2821_1), .Y(N2821) );
  AND2X1 gate833_1 ( .A(N898), .B(N283), .Y(N2824_1) );
  AND2X1 gate833 ( .A(N2789), .B(N2824_1), .Y(N2824) );
  NAND2X1 gate834 ( .A(N1965), .B(N2808), .Y(N2827) );
  NAND2X1 gate835 ( .A(N1968), .B(N2810), .Y(N2828) );
  AND2X1 gate836_1 ( .A(N79), .B(N283), .Y(N2829_1) );
  AND2X1 gate836 ( .A(N2789), .B(N2829_1), .Y(N2829) );
  NAND2X1 gate837 ( .A(N2807), .B(N2827), .Y(N2843) );
  NAND2X1 gate838 ( .A(N2809), .B(N2828), .Y(N2846) );
  NAND2X1 gate839 ( .A(N2812), .B(N2076), .Y(N2850) );
  NAND2X1 gate840 ( .A(N2815), .B(N2077), .Y(N2851) );
  NAND2X1 gate841 ( .A(N2818), .B(N1915), .Y(N2852) );
  NAND2X1 gate842 ( .A(N2821), .B(N1857), .Y(N2853) );
  NAND2X1 gate843 ( .A(N2824), .B(N1938), .Y(N2854) );
  INVX1 gate844 ( .A(N2812), .Y(N2857) );
  INVX1 gate845 ( .A(N2815), .Y(N2858) );
  INVX1 gate846 ( .A(N2818), .Y(N2859) );
  INVX1 gate847 ( .A(N2821), .Y(N2860) );
  INVX1 gate848 ( .A(N2824), .Y(N2861) );
  INVX1 gate849 ( .A(N2829), .Y(N2862) );
  NAND2X1 gate850 ( .A(N2829), .B(N1985), .Y(N2863) );
  NAND2X1 gate851 ( .A(N2052), .B(N2857), .Y(N2866) );
  NAND2X1 gate852 ( .A(N2055), .B(N2858), .Y(N2867) );
  NAND2X1 gate853 ( .A(N1866), .B(N2859), .Y(N2868) );
  NAND2X1 gate854 ( .A(N1818), .B(N2860), .Y(N2869) );
  NAND2X1 gate855 ( .A(N1902), .B(N2861), .Y(N2870) );
  NAND2X1 gate856 ( .A(N2843), .B(N886), .Y(N2871) );
  INVX1 gate857 ( .A(N2843), .Y(N2872) );
  NAND2X1 gate858 ( .A(N2846), .B(N887), .Y(N2873) );
  INVX1 gate859 ( .A(N2846), .Y(N2874) );
  NAND2X1 gate860 ( .A(N1933), .B(N2862), .Y(N2875) );
  NAND2X1 gate861 ( .A(N2866), .B(N2850), .Y(N2876) );
  NAND2X1 gate862 ( .A(N2867), .B(N2851), .Y(N2877) );
  NAND2X1 gate863 ( .A(N2868), .B(N2852), .Y(N2878) );
  NAND2X1 gate864 ( .A(N2869), .B(N2853), .Y(N2879) );
  NAND2X1 gate865 ( .A(N2870), .B(N2854), .Y(N2880) );
  NAND2X1 gate866 ( .A(N682), .B(N2872), .Y(N2881) );
  NAND2X1 gate867 ( .A(N685), .B(N2874), .Y(N2882) );
  NAND2X1 gate868 ( .A(N2875), .B(N2863), .Y(N2883) );
  AND2X1 gate869 ( .A(N2876), .B(N550), .Y(N2886) );
  AND2X1 gate870 ( .A(N551), .B(N2877), .Y(N2887) );
  AND2X1 gate871 ( .A(N553), .B(N2878), .Y(N2888) );
  AND2X1 gate872 ( .A(N2879), .B(N554), .Y(N2889) );
  AND2X1 gate873 ( .A(N555), .B(N2880), .Y(N2890) );
  NAND2X1 gate874 ( .A(N2871), .B(N2881), .Y(N2891) );
  NAND2X1 gate875 ( .A(N2873), .B(N2882), .Y(N2892) );
  NAND2X1 gate876 ( .A(N2883), .B(N1461), .Y(N2895) );
  INVX1 gate877 ( .A(N2883), .Y(N2896) );
  NAND2X1 gate878 ( .A(N1383), .B(N2896), .Y(N2897) );
  NAND2X1 gate879 ( .A(N2895), .B(N2897), .Y(N2898) );
  AND2X1 gate880 ( .A(N2898), .B(N552), .Y(N2899) );
endmodule


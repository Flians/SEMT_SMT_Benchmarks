
module c3540_synth ( N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, 
        N107, N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, 
        N190, N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, 
        N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, 
        N349, N350, N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, 
        N4667, N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, 
        N5192, N5231, N5360, N5361 );
  input N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116,
         N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190,
         N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264,
         N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330,
         N343, N349, N350;
  output N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815,
         N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231,
         N5360, N5361;
  wire   N655, N665, N670, N679, N683, N686, N690, N699, N702, N706, N715,
         N724, N727, N736, N740, N749, N753, N763, N768, N769, N772, N779,
         N782, N786, N793, N794, N798, N803, N820, N821, N825, N829, N832,
         N835, N836, N839, N842, N845, N848, N851, N854, N858, N861, N864,
         N867, N870, N874, N877, N880, N883, N886, N889, N890, N891, N892,
         N895, N896, N913, N914, N915, N916, N917, N920, N923, N926, N929,
         N932, N935, N938, N941, N944, N947, N950, N953, N956, N959, N962,
         N965, N1067, N1117, N1179, N1196, N1197, N1202, N1219, N1250, N1251,
         N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261,
         N1262, N1263, N1264, N1267, N1268, N1271, N1272, N1273, N1276, N1279,
         N1298, N1302, N1306, N1315, N1322, N1325, N1328, N1331, N1334, N1337,
         N1338, N1339, N1340, N1343, N1344, N1345, N1346, N1347, N1348, N1349,
         N1350, N1351, N1352, N1353, N1358, N1363, N1366, N1369, N1384, N1401,
         N1402, N1403, N1404, N1405, N1406, N1407, N1408, N1409, N1426, N1427,
         N1452, N1459, N1460, N1461, N1464, N1467, N1468, N1469, N1470, N1471,
         N1474, N1475, N1478, N1481, N1484, N1487, N1490, N1493, N1496, N1499,
         N1502, N1505, N1507, N1508, N1509, N1510, N1511, N1512, N1520, N1562,
         N1579, N1580, N1581, N1582, N1583, N1584, N1585, N1586, N1587, N1588,
         N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598,
         N1599, N1600, N1643, N1644, N1645, N1646, N1647, N1648, N1649, N1650,
         N1667, N1670, N1673, N1674, N1675, N1676, N1677, N1678, N1679, N1680,
         N1691, N1692, N1693, N1694, N1714, N1715, N1718, N1721, N1722, N1725,
         N1726, N1727, N1728, N1729, N1730, N1731, N1735, N1736, N1737, N1738,
         N1747, N1756, N1761, N1764, N1765, N1766, N1767, N1768, N1769, N1770,
         N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794, N1795, N1796,
         N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1806, N1809, N1812,
         N1815, N1818, N1821, N1824, N1833, N1842, N1843, N1844, N1845, N1846,
         N1847, N1848, N1849, N1850, N1851, N1852, N1853, N1854, N1855, N1856,
         N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864, N1869, N1870,
         N1873, N1874, N1875, N1878, N1879, N1880, N1883, N1884, N1885, N1888,
         N1889, N1890, N1893, N1894, N1895, N1898, N1899, N1900, N1903, N1904,
         N1905, N1908, N1909, N1912, N1913, N1917, N1922, N1926, N1930, N1933,
         N1936, N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1960,
         N1961, N1966, N1981, N1982, N1983, N1986, N1987, N1988, N1989, N1990,
         N1991, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030,
         N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, N2043, N2052,
         N2057, N2068, N2073, N2078, N2083, N2088, N2093, N2098, N2103, N2121,
         N2122, N2123, N2124, N2125, N2126, N2127, N2128, N2133, N2134, N2135,
         N2136, N2137, N2138, N2139, N2141, N2142, N2143, N2144, N2145, N2146,
         N2147, N2148, N2149, N2150, N2151, N2152, N2153, N2154, N2155, N2156,
         N2157, N2158, N2175, N2178, N2179, N2180, N2181, N2183, N2184, N2185,
         N2188, N2191, N2194, N2197, N2200, N2203, N2206, N2209, N2210, N2211,
         N2212, N2221, N2230, N2231, N2232, N2233, N2234, N2235, N2236, N2237,
         N2238, N2239, N2240, N2241, N2242, N2243, N2244, N2245, N2270, N2277,
         N2282, N2287, N2294, N2299, N2304, N2307, N2310, N2313, N2316, N2319,
         N2322, N2325, N2328, N2331, N2334, N2341, N2342, N2347, N2348, N2349,
         N2350, N2351, N2352, N2353, N2354, N2355, N2374, N2375, N2376, N2379,
         N2398, N2417, N2418, N2419, N2420, N2421, N2422, N2425, N2426, N2427,
         N2430, N2431, N2432, N2435, N2436, N2437, N2438, N2439, N2440, N2443,
         N2444, N2445, N2448, N2449, N2450, N2467, N2468, N2469, N2470, N2471,
         N2474, N2475, N2476, N2477, N2478, N2481, N2482, N2483, N2486, N2487,
         N2488, N2497, N2506, N2515, N2524, N2533, N2542, N2551, N2560, N2569,
         N2578, N2587, N2596, N2605, N2614, N2623, N2632, N2633, N2634, N2635,
         N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645,
         N2646, N2647, N2648, N2652, N2656, N2659, N2662, N2666, N2670, N2673,
         N2677, N2681, N2684, N2688, N2692, N2697, N2702, N2706, N2710, N2715,
         N2719, N2723, N2728, N2729, N2730, N2731, N2732, N2733, N2734, N2735,
         N2736, N2737, N2738, N2739, N2740, N2741, N2742, N2743, N2744, N2745,
         N2746, N2748, N2749, N2750, N2751, N2754, N2755, N2756, N2757, N2758,
         N2761, N2764, N2768, N2769, N2898, N2899, N2900, N2901, N2962, N2966,
         N2967, N2970, N2973, N2977, N2980, N2984, N2985, N2986, N2987, N2988,
         N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998,
         N2999, N3000, N3001, N3002, N3003, N3004, N3005, N3006, N3007, N3008,
         N3009, N3010, N3011, N3012, N3013, N3014, N3015, N3016, N3017, N3018,
         N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028,
         N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3036, N3037, N3038,
         N3039, N3040, N3041, N3042, N3043, N3044, N3045, N3046, N3047, N3048,
         N3049, N3050, N3051, N3052, N3053, N3054, N3055, N3056, N3057, N3058,
         N3059, N3060, N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068,
         N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078,
         N3079, N3080, N3081, N3082, N3083, N3084, N3085, N3086, N3087, N3088,
         N3089, N3090, N3091, N3092, N3093, N3094, N3095, N3096, N3097, N3098,
         N3099, N3100, N3101, N3102, N3103, N3104, N3105, N3106, N3107, N3108,
         N3109, N3110, N3111, N3112, N3115, N3118, N3119, N3122, N3125, N3128,
         N3131, N3134, N3135, N3138, N3141, N3142, N3145, N3148, N3149, N3152,
         N3155, N3158, N3161, N3164, N3165, N3168, N3171, N3172, N3175, N3178,
         N3181, N3184, N3187, N3190, N3191, N3192, N3193, N3194, N3196, N3206,
         N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3216,
         N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224, N3225, N3226,
         N3227, N3228, N3229, N3230, N3231, N3232, N3233, N3234, N3235, N3236,
         N3237, N3238, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246,
         N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254, N3255, N3256,
         N3257, N3258, N3259, N3260, N3261, N3262, N3263, N3264, N3265, N3266,
         N3267, N3268, N3269, N3270, N3271, N3272, N3273, N3274, N3275, N3276,
         N3277, N3278, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286,
         N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294, N3295, N3296,
         N3297, N3298, N3299, N3300, N3301, N3302, N3303, N3304, N3305, N3306,
         N3307, N3308, N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316,
         N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326,
         N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3383, N3384,
         N3387, N3388, N3389, N3390, N3391, N3392, N3393, N3394, N3395, N3396,
         N3397, N3398, N3399, N3400, N3401, N3402, N3403, N3404, N3405, N3406,
         N3407, N3410, N3413, N3414, N3415, N3419, N3423, N3426, N3429, N3430,
         N3431, N3434, N3437, N3438, N3439, N3442, N3445, N3446, N3447, N3451,
         N3455, N3458, N3461, N3462, N3463, N3466, N3469, N3470, N3471, N3472,
         N3475, N3478, N3481, N3484, N3487, N3490, N3493, N3496, N3499, N3502,
         N3505, N3508, N3511, N3514, N3517, N3520, N3523, N3534, N3535, N3536,
         N3537, N3538, N3539, N3540, N3541, N3542, N3543, N3544, N3545, N3546,
         N3547, N3548, N3549, N3550, N3551, N3552, N3557, N3568, N3573, N3578,
         N3589, N3594, N3605, N3626, N3627, N3628, N3629, N3630, N3631, N3632,
         N3633, N3634, N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642,
         N3643, N3644, N3645, N3648, N3651, N3652, N3653, N3654, N3657, N3658,
         N3661, N3662, N3663, N3664, N3667, N3670, N3671, N3672, N3673, N3676,
         N3677, N3680, N3681, N3682, N3685, N3686, N3687, N3688, N3689, N3690,
         N3693, N3694, N3695, N3696, N3697, N3700, N3703, N3704, N3705, N3706,
         N3707, N3708, N3711, N3712, N3713, N3714, N3715, N3716, N3717, N3718,
         N3719, N3720, N3721, N3731, N3734, N3740, N3743, N3753, N3756, N3762,
         N3765, N3766, N3773, N3774, N3775, N3776, N3777, N3778, N3779, N3780,
         N3786, N3789, N3800, N3803, N3809, N3812, N3815, N3818, N3821, N3824,
         N3827, N3830, N3834, N3835, N3838, N3845, N3850, N3855, N3858, N3861,
         N3865, N3868, N3884, N3885, N3894, N3895, N3898, N3899, N3906, N3911,
         N3912, N3913, N3916, N3917, N3920, N3921, N3924, N3925, N3926, N3930,
         N3931, N3932, N3935, N3936, N3937, N3940, N3947, N3948, N3950, N3953,
         N3956, N3959, N3962, N3965, N3968, N3971, N3974, N3977, N3980, N3983,
         N3992, N3996, N4013, N4029, N4030, N4031, N4032, N4033, N4034, N4035,
         N4042, N4043, N4044, N4045, N4046, N4047, N4048, N4049, N4050, N4051,
         N4052, N4053, N4054, N4055, N4056, N4057, N4058, N4059, N4062, N4065,
         N4066, N4067, N4070, N4073, N4074, N4075, N4076, N4077, N4078, N4079,
         N4080, N4085, N4086, N4088, N4090, N4091, N4094, N4098, N4101, N4104,
         N4105, N4106, N4107, N4108, N4109, N4110, N4111, N4112, N4113, N4114,
         N4115, N4116, N4119, N4122, N4123, N4126, N4127, N4128, N4139, N4142,
         N4146, N4147, N4148, N4149, N4150, N4151, N4152, N4153, N4154, N4161,
         N4167, N4174, N4182, N4186, N4189, N4190, N4191, N4192, N4193, N4194,
         N4195, N4196, N4197, N4200, N4203, N4209, N4213, N4218, N4223, N4238,
         N4239, N4241, N4242, N4247, N4251, N4252, N4253, N4254, N4255, N4256,
         N4257, N4258, N4283, N4284, N4287, N4291, N4295, N4296, N4299, N4303,
         N4304, N4305, N4310, N4316, N4317, N4318, N4319, N4322, N4325, N4326,
         N4327, N4328, N4329, N4330, N4331, N4335, N4338, N4341, N4344, N4347,
         N4350, N4353, N4356, N4359, N4362, N4365, N4368, N4371, N4376, N4377,
         N4387, N4390, N4393, N4398, N4413, N4416, N4421, N4427, N4430, N4435,
         N4442, N4443, N4446, N4447, N4448, N4452, N4458, N4461, N4462, N4463,
         N4464, N4465, N4468, N4472, N4475, N4479, N4484, N4486, N4487, N4491,
         N4493, N4496, N4497, N4498, N4503, N4506, N4507, N4508, N4509, N4510,
         N4511, N4515, N4526, N4527, N4528, N4529, N4530, N4531, N4534, N4537,
         N4540, N4545, N4549, N4552, N4555, N4558, N4559, N4562, N4563, N4564,
         N4568, N4569, N4572, N4573, N4576, N4581, N4584, N4587, N4588, N4593,
         N4596, N4597, N4599, N4602, N4603, N4608, N4613, N4616, N4619, N4623,
         N4628, N4629, N4630, N4635, N4636, N4640, N4641, N4642, N4643, N4644,
         N4647, N4650, N4656, N4659, N4664, N4668, N4669, N4670, N4673, N4674,
         N4675, N4676, N4677, N4678, N4679, N4687, N4688, N4691, N4694, N4697,
         N4700, N4704, N4705, N4706, N4707, N4708, N4711, N4716, N4717, N4721,
         N4722, N4726, N4727, N4730, N4733, N4740, N4743, N4747, N4748, N4749,
         N4750, N4753, N4754, N4755, N4756, N4757, N4769, N4772, N4775, N4778,
         N4786, N4787, N4788, N4789, N4794, N4797, N4800, N4805, N4808, N4812,
         N4816, N4817, N4818, N4822, N4823, N4826, N4829, N4830, N4831, N4838,
         N4844, N4847, N4850, N4854, N4859, N4860, N4868, N4870, N4872, N4873,
         N4876, N4880, N4885, N4889, N4895, N4896, N4897, N4898, N4899, N4900,
         N4901, N4902, N4904, N4905, N4906, N4907, N4913, N4916, N4920, N4921,
         N4924, N4925, N4926, N4928, N4929, N4930, N4931, N4937, N4940, N4946,
         N4949, N4950, N4951, N4952, N4953, N4954, N4957, N4964, N4965, N4968,
         N4969, N4970, N4973, N4978, N4979, N4980, N4981, N4982, N4983, N4984,
         N4985, N4988, N4991, N4996, N4999, N5007, N5010, N5013, N5018, N5021,
         N5026, N5029, N5030, N5039, N5042, N5046, N5050, N5055, N5058, N5061,
         N5066, N5070, N5080, N5085, N5094, N5095, N5097, N5103, N5108, N5109,
         N5110, N5111, N5114, N5117, N5122, N5125, N5128, N5133, N5136, N5139,
         N5145, N5151, N5154, N5159, N5160, N5163, N5166, N5173, N5174, N5177,
         N5182, N5183, N5184, N5188, N5193, N5196, N5197, N5198, N5199, N5201,
         N5203, N5205, N5209, N5212, N5215, N5217, N5219, N5220, N5221, N5222,
         N5223, N5224, N5225, N5228, N5232, N5233, N5234, N5235, N5236, N5240,
         N5242, N5243, N5245, N5246, N5250, N5253, N5254, N5257, N5258, N5261,
         N5266, N5269, N5277, N5278, N5279, N5283, N5284, N5285, N5286, N5289,
         N5292, N5295, N5298, N5303, N5306, N5309, N5312, N5313, N5322, N5323,
         N5324, N5327, N5332, N5335, N5340, N5341, N5344, N5345, N5348, N5349,
         N5350, N5351, N5352, N5353, N5354, N5355, N5356, N5357, N5358, N5359,
         N1250_1, N1315_1, N1325_1, N1340_1, N1452_1, N1507_1, N1507_2,
         N1508_1, N1508_2, N1667_1, N1670_1, N1761_1, N1761_2, N1913_1,
         N1922_1, N1986_1, N1987_1, N1988_1, N1989_1, N1990_1, N1991_1,
         N2068_1, N2073_1, N2078_1, N2083_1, N2088_1, N2093_1, N2098_1,
         N2103_1, N2148_1, N2148_2, N2238_1, N2239_1, N2240_1, N2241_1,
         N2242_1, N2243_1, N2244_1, N2245_1, N2348_1, N2417_1, N2418_1,
         N2420_1, N2421_1, N2425_1, N2426_1, N2430_1, N2431_1, N2435_1,
         N2436_1, N2438_1, N2439_1, N2443_1, N2444_1, N2448_1, N2449_1,
         N2648_1, N2656_1, N2659_1, N2662_1, N2670_1, N2673_1, N2681_1,
         N2684_1, N2692_1, N2697_1, N2702_1, N2710_1, N2715_1, N2723_1,
         N2745_1, N2768_1, N2769_1, N3194_1, N3194_2, N3194_3, N3206_1,
         N3383_1, N3383_2, N3383_3, N3390_1, N3390_2, N3390_3, N3391_1,
         N3391_2, N3391_3, N3392_1, N3392_2, N3392_3, N3393_1, N3393_2,
         N3393_3, N3394_1, N3394_2, N3394_3, N3395_1, N3395_2, N3395_3,
         N3396_1, N3396_2, N3396_3, N3397_1, N3397_2, N3397_3, N3398_1,
         N3398_2, N3398_3, N3399_1, N3399_2, N3399_3, N3400_1, N3400_2,
         N3400_3, N3401_1, N3401_2, N3401_3, N3402_1, N3402_2, N3402_3,
         N3403_1, N3403_2, N3403_3, N3404_1, N3404_2, N3404_3, N3405_1,
         N3405_2, N3405_3, N3407_1, N3410_1, N3413_1, N3414_1, N3415_1,
         N3423_1, N3426_1, N3429_1, N3430_1, N3431_1, N3434_1, N3437_1,
         N3438_1, N3439_1, N3442_1, N3445_1, N3446_1, N3447_1, N3455_1,
         N3458_1, N3461_1, N3462_1, N3463_1, N3466_1, N3469_1, N3470_1,
         N3535_1, N3557_1, N3568_1, N3573_1, N3578_1, N3589_1, N3594_1,
         N3634_1, N3645_1, N3648_1, N3651_1, N3652_1, N3664_1, N3667_1,
         N3670_1, N3671_1, N3711_1, N3712_1, N3731_1, N3753_1, N3926_1,
         N3926_2, N3931_1, N3931_2, N3932_1, N3932_2, N3936_1, N3936_2,
         N3992_1, N3992_2, N3996_1, N3996_2, N4316_1, N4318_1, N4331_1,
         N4443_1, N4443_2, N4448_1, N4448_2, N4503_1, N4503_2, N4545_1,
         N4587_1, N4608_1, N4727_1, N4876_1, N4901_1, N4901_2, N4964_1,
         N4982_1, N4982_2, N4988_1, N4996_1, N5018_1, N5050_1, N5058_1,
         N5066_1, N5066_2, N5080_1, N5133_1, N5133_2, N5136_1, N5277_1,
         N5278_1, N5285_1, N5286_1, N5298_1, N5298_2;

  BUFX2 gate1 ( .A(N50), .Y(N655) );
  INVX1 gate2 ( .A(N50), .Y(N665) );
  BUFX2 gate3 ( .A(N58), .Y(N670) );
  INVX1 gate4 ( .A(N58), .Y(N679) );
  BUFX2 gate5 ( .A(N68), .Y(N683) );
  INVX1 gate6 ( .A(N68), .Y(N686) );
  BUFX2 gate7 ( .A(N68), .Y(N690) );
  BUFX2 gate8 ( .A(N77), .Y(N699) );
  INVX1 gate9 ( .A(N77), .Y(N702) );
  BUFX2 gate10 ( .A(N77), .Y(N706) );
  BUFX2 gate11 ( .A(N87), .Y(N715) );
  INVX1 gate12 ( .A(N87), .Y(N724) );
  BUFX2 gate13 ( .A(N97), .Y(N727) );
  INVX1 gate14 ( .A(N97), .Y(N736) );
  BUFX2 gate15 ( .A(N107), .Y(N740) );
  INVX1 gate16 ( .A(N107), .Y(N749) );
  BUFX2 gate17 ( .A(N116), .Y(N753) );
  INVX1 gate18 ( .A(N116), .Y(N763) );
  OR2X1 gate19 ( .A(N257), .B(N264), .Y(N768) );
  INVX1 gate20 ( .A(N1), .Y(N769) );
  BUFX2 gate21 ( .A(N1), .Y(N772) );
  INVX1 gate22 ( .A(N1), .Y(N779) );
  BUFX2 gate23 ( .A(N13), .Y(N782) );
  INVX1 gate24 ( .A(N13), .Y(N786) );
  AND2X1 gate25 ( .A(N13), .B(N20), .Y(N793) );
  INVX1 gate26 ( .A(N20), .Y(N794) );
  BUFX2 gate27 ( .A(N20), .Y(N798) );
  INVX1 gate28 ( .A(N20), .Y(N803) );
  INVX1 gate29 ( .A(N33), .Y(N820) );
  BUFX2 gate30 ( .A(N33), .Y(N821) );
  INVX1 gate31 ( .A(N33), .Y(N825) );
  AND2X1 gate32 ( .A(N33), .B(N41), .Y(N829) );
  INVX1 gate33 ( .A(N41), .Y(N832) );
  OR2X1 gate34 ( .A(N41), .B(N45), .Y(N835) );
  BUFX2 gate35 ( .A(N45), .Y(N836) );
  INVX1 gate36 ( .A(N45), .Y(N839) );
  INVX1 gate37 ( .A(N50), .Y(N842) );
  BUFX2 gate38 ( .A(N58), .Y(N845) );
  INVX1 gate39 ( .A(N58), .Y(N848) );
  BUFX2 gate40 ( .A(N68), .Y(N851) );
  INVX1 gate41 ( .A(N68), .Y(N854) );
  BUFX2 gate42 ( .A(N87), .Y(N858) );
  INVX1 gate43 ( .A(N87), .Y(N861) );
  BUFX2 gate44 ( .A(N97), .Y(N864) );
  INVX1 gate45 ( .A(N97), .Y(N867) );
  INVX1 gate46 ( .A(N107), .Y(N870) );
  BUFX2 gate47 ( .A(N1), .Y(N874) );
  BUFX2 gate48 ( .A(N68), .Y(N877) );
  BUFX2 gate49 ( .A(N107), .Y(N880) );
  INVX1 gate50 ( .A(N20), .Y(N883) );
  BUFX2 gate51 ( .A(N190), .Y(N886) );
  INVX1 gate52 ( .A(N200), .Y(N889) );
  AND2X1 gate53 ( .A(N20), .B(N200), .Y(N890) );
  NAND2X1 gate54 ( .A(N20), .B(N200), .Y(N891) );
  AND2X1 gate55 ( .A(N20), .B(N179), .Y(N892) );
  INVX1 gate56 ( .A(N20), .Y(N895) );
  OR2X1 gate57 ( .A(N349), .B(N33), .Y(N896) );
  NAND2X1 gate58 ( .A(N1), .B(N13), .Y(N913) );
  NAND3X1 gate59 ( .A(N1), .B(N20), .C(N33), .Y(N914) );
  INVX1 gate60 ( .A(N20), .Y(N915) );
  INVX1 gate61 ( .A(N33), .Y(N916) );
  BUFX2 gate62 ( .A(N179), .Y(N917) );
  INVX1 gate63 ( .A(N213), .Y(N920) );
  BUFX2 gate64 ( .A(N343), .Y(N923) );
  BUFX2 gate65 ( .A(N226), .Y(N926) );
  BUFX2 gate66 ( .A(N232), .Y(N929) );
  BUFX2 gate67 ( .A(N238), .Y(N932) );
  BUFX2 gate68 ( .A(N244), .Y(N935) );
  BUFX2 gate69 ( .A(N250), .Y(N938) );
  BUFX2 gate70 ( .A(N257), .Y(N941) );
  BUFX2 gate71 ( .A(N264), .Y(N944) );
  BUFX2 gate72 ( .A(N270), .Y(N947) );
  BUFX2 gate73 ( .A(N50), .Y(N950) );
  BUFX2 gate74 ( .A(N58), .Y(N953) );
  BUFX2 gate75 ( .A(N58), .Y(N956) );
  BUFX2 gate76 ( .A(N97), .Y(N959) );
  BUFX2 gate77 ( .A(N97), .Y(N962) );
  BUFX2 gate78 ( .A(N330), .Y(N965) );
  AND2X1 gate79 ( .A(N250), .B(N768), .Y(N1067) );
  OR2X1 gate80 ( .A(N820), .B(N20), .Y(N1117) );
  OR2X1 gate81 ( .A(N895), .B(N169), .Y(N1179) );
  INVX1 gate82 ( .A(N793), .Y(N1196) );
  OR2X1 gate83 ( .A(N915), .B(N1), .Y(N1197) );
  AND2X1 gate84 ( .A(N913), .B(N914), .Y(N1202) );
  OR2X1 gate85 ( .A(N916), .B(N1), .Y(N1219) );
  AND2X1 gate86_1 ( .A(N842), .B(N848), .Y(N1250_1) );
  AND2X1 gate86 ( .A(N854), .B(N1250_1), .Y(N1250) );
  NAND2X1 gate87 ( .A(N226), .B(N655), .Y(N1251) );
  NAND2X1 gate88 ( .A(N232), .B(N670), .Y(N1252) );
  NAND2X1 gate89 ( .A(N238), .B(N690), .Y(N1253) );
  NAND2X1 gate90 ( .A(N244), .B(N706), .Y(N1254) );
  NAND2X1 gate91 ( .A(N250), .B(N715), .Y(N1255) );
  NAND2X1 gate92 ( .A(N257), .B(N727), .Y(N1256) );
  NAND2X1 gate93 ( .A(N264), .B(N740), .Y(N1257) );
  NAND2X1 gate94 ( .A(N270), .B(N753), .Y(N1258) );
  INVX1 gate95 ( .A(N926), .Y(N1259) );
  INVX1 gate96 ( .A(N929), .Y(N1260) );
  INVX1 gate97 ( .A(N932), .Y(N1261) );
  INVX1 gate98 ( .A(N935), .Y(N1262) );
  NAND2X1 gate99 ( .A(N679), .B(N686), .Y(N1263) );
  NAND2X1 gate100 ( .A(N736), .B(N749), .Y(N1264) );
  NAND2X1 gate101 ( .A(N683), .B(N699), .Y(N1267) );
  BUFX2 gate102 ( .A(N665), .Y(N1268) );
  INVX1 gate103 ( .A(N953), .Y(N1271) );
  INVX1 gate104 ( .A(N959), .Y(N1272) );
  BUFX2 gate105 ( .A(N839), .Y(N1273) );
  BUFX2 gate106 ( .A(N839), .Y(N1276) );
  BUFX2 gate107 ( .A(N782), .Y(N1279) );
  BUFX2 gate108 ( .A(N825), .Y(N1298) );
  BUFX2 gate109 ( .A(N832), .Y(N1302) );
  AND2X1 gate110 ( .A(N779), .B(N835), .Y(N1306) );
  AND2X1 gate111_1 ( .A(N779), .B(N836), .Y(N1315_1) );
  AND2X1 gate111 ( .A(N832), .B(N1315_1), .Y(N1315) );
  AND2X1 gate112 ( .A(N769), .B(N836), .Y(N1322) );
  AND2X1 gate113_1 ( .A(N772), .B(N786), .Y(N1325_1) );
  AND2X1 gate113 ( .A(N798), .B(N1325_1), .Y(N1325) );
  NAND3X1 gate114 ( .A(N772), .B(N786), .C(N798), .Y(N1328) );
  NAND2X1 gate115 ( .A(N772), .B(N786), .Y(N1331) );
  BUFX2 gate116 ( .A(N874), .Y(N1334) );
  NAND3X1 gate117 ( .A(N782), .B(N794), .C(N45), .Y(N1337) );
  NAND3X1 gate118 ( .A(N842), .B(N848), .C(N854), .Y(N1338) );
  INVX1 gate119 ( .A(N956), .Y(N1339) );
  AND2X1 gate120_1 ( .A(N861), .B(N867), .Y(N1340_1) );
  AND2X1 gate120 ( .A(N870), .B(N1340_1), .Y(N1340) );
  NAND3X1 gate121 ( .A(N861), .B(N867), .C(N870), .Y(N1343) );
  INVX1 gate122 ( .A(N962), .Y(N1344) );
  INVX1 gate123 ( .A(N803), .Y(N1345) );
  INVX1 gate124 ( .A(N803), .Y(N1346) );
  INVX1 gate125 ( .A(N803), .Y(N1347) );
  INVX1 gate126 ( .A(N803), .Y(N1348) );
  INVX1 gate127 ( .A(N803), .Y(N1349) );
  INVX1 gate128 ( .A(N803), .Y(N1350) );
  INVX1 gate129 ( .A(N803), .Y(N1351) );
  INVX1 gate130 ( .A(N803), .Y(N1352) );
  OR2X1 gate131 ( .A(N883), .B(N886), .Y(N1353) );
  NOR2X1 gate132 ( .A(N883), .B(N886), .Y(N1358) );
  BUFX2 gate133 ( .A(N892), .Y(N1363) );
  INVX1 gate134 ( .A(N892), .Y(N1366) );
  BUFX2 gate135 ( .A(N821), .Y(N1369) );
  BUFX2 gate136 ( .A(N825), .Y(N1384) );
  INVX1 gate137 ( .A(N896), .Y(N1401) );
  INVX1 gate138 ( .A(N896), .Y(N1402) );
  INVX1 gate139 ( .A(N896), .Y(N1403) );
  INVX1 gate140 ( .A(N896), .Y(N1404) );
  INVX1 gate141 ( .A(N896), .Y(N1405) );
  INVX1 gate142 ( .A(N896), .Y(N1406) );
  INVX1 gate143 ( .A(N896), .Y(N1407) );
  INVX1 gate144 ( .A(N896), .Y(N1408) );
  OR2X1 gate145 ( .A(N1), .B(N1196), .Y(N1409) );
  INVX1 gate146 ( .A(N829), .Y(N1426) );
  INVX1 gate147 ( .A(N829), .Y(N1427) );
  AND2X1 gate148_1 ( .A(N769), .B(N782), .Y(N1452_1) );
  AND2X1 gate148 ( .A(N794), .B(N1452_1), .Y(N1452) );
  INVX1 gate149 ( .A(N917), .Y(N1459) );
  INVX1 gate150 ( .A(N965), .Y(N1460) );
  OR2X1 gate151 ( .A(N920), .B(N923), .Y(N1461) );
  NOR2X1 gate152 ( .A(N920), .B(N923), .Y(N1464) );
  INVX1 gate153 ( .A(N938), .Y(N1467) );
  INVX1 gate154 ( .A(N941), .Y(N1468) );
  INVX1 gate155 ( .A(N944), .Y(N1469) );
  INVX1 gate156 ( .A(N947), .Y(N1470) );
  BUFX2 gate157 ( .A(N679), .Y(N1471) );
  INVX1 gate158 ( .A(N950), .Y(N1474) );
  BUFX2 gate159 ( .A(N686), .Y(N1475) );
  BUFX2 gate160 ( .A(N702), .Y(N1478) );
  BUFX2 gate161 ( .A(N724), .Y(N1481) );
  BUFX2 gate162 ( .A(N736), .Y(N1484) );
  BUFX2 gate163 ( .A(N749), .Y(N1487) );
  BUFX2 gate164 ( .A(N763), .Y(N1490) );
  BUFX2 gate165 ( .A(N877), .Y(N1493) );
  BUFX2 gate166 ( .A(N877), .Y(N1496) );
  BUFX2 gate167 ( .A(N880), .Y(N1499) );
  BUFX2 gate168 ( .A(N880), .Y(N1502) );
  NAND2X1 gate169 ( .A(N702), .B(N1250), .Y(N1505) );
  AND2X1 gate170_1 ( .A(N1251), .B(N1252), .Y(N1507_1) );
  AND2X1 gate170_2 ( .A(N1253), .B(N1254), .Y(N1507_2) );
  AND2X1 gate170 ( .A(N1507_1), .B(N1507_2), .Y(N1507) );
  AND2X1 gate171_1 ( .A(N1255), .B(N1256), .Y(N1508_1) );
  AND2X1 gate171_2 ( .A(N1257), .B(N1258), .Y(N1508_2) );
  AND2X1 gate171 ( .A(N1508_1), .B(N1508_2), .Y(N1508) );
  NAND2X1 gate172 ( .A(N929), .B(N1259), .Y(N1509) );
  NAND2X1 gate173 ( .A(N926), .B(N1260), .Y(N1510) );
  NAND2X1 gate174 ( .A(N935), .B(N1261), .Y(N1511) );
  NAND2X1 gate175 ( .A(N932), .B(N1262), .Y(N1512) );
  AND2X1 gate176 ( .A(N655), .B(N1263), .Y(N1520) );
  AND2X1 gate177 ( .A(N874), .B(N1337), .Y(N1562) );
  INVX1 gate178 ( .A(N1117), .Y(N1579) );
  AND2X1 gate179 ( .A(N803), .B(N1117), .Y(N1580) );
  AND2X1 gate180 ( .A(N1338), .B(N1345), .Y(N1581) );
  INVX1 gate181 ( .A(N1117), .Y(N1582) );
  AND2X1 gate182 ( .A(N803), .B(N1117), .Y(N1583) );
  INVX1 gate183 ( .A(N1117), .Y(N1584) );
  AND2X1 gate184 ( .A(N803), .B(N1117), .Y(N1585) );
  AND2X1 gate185 ( .A(N854), .B(N1347), .Y(N1586) );
  INVX1 gate186 ( .A(N1117), .Y(N1587) );
  AND2X1 gate187 ( .A(N803), .B(N1117), .Y(N1588) );
  AND2X1 gate188 ( .A(N77), .B(N1348), .Y(N1589) );
  INVX1 gate189 ( .A(N1117), .Y(N1590) );
  AND2X1 gate190 ( .A(N803), .B(N1117), .Y(N1591) );
  AND2X1 gate191 ( .A(N1343), .B(N1349), .Y(N1592) );
  INVX1 gate192 ( .A(N1117), .Y(N1593) );
  AND2X1 gate193 ( .A(N803), .B(N1117), .Y(N1594) );
  INVX1 gate194 ( .A(N1117), .Y(N1595) );
  AND2X1 gate195 ( .A(N803), .B(N1117), .Y(N1596) );
  AND2X1 gate196 ( .A(N870), .B(N1351), .Y(N1597) );
  INVX1 gate197 ( .A(N1117), .Y(N1598) );
  AND2X1 gate198 ( .A(N803), .B(N1117), .Y(N1599) );
  AND2X1 gate199 ( .A(N116), .B(N1352), .Y(N1600) );
  AND2X1 gate200 ( .A(N222), .B(N1401), .Y(N1643) );
  AND2X1 gate201 ( .A(N223), .B(N1402), .Y(N1644) );
  AND2X1 gate202 ( .A(N226), .B(N1403), .Y(N1645) );
  AND2X1 gate203 ( .A(N232), .B(N1404), .Y(N1646) );
  AND2X1 gate204 ( .A(N238), .B(N1405), .Y(N1647) );
  AND2X1 gate205 ( .A(N244), .B(N1406), .Y(N1648) );
  AND2X1 gate206 ( .A(N250), .B(N1407), .Y(N1649) );
  AND2X1 gate207 ( .A(N257), .B(N1408), .Y(N1650) );
  AND2X1 gate208_1 ( .A(N1), .B(N13), .Y(N1667_1) );
  AND2X1 gate208 ( .A(N1426), .B(N1667_1), .Y(N1667) );
  AND2X1 gate209_1 ( .A(N1), .B(N13), .Y(N1670_1) );
  AND2X1 gate209 ( .A(N1427), .B(N1670_1), .Y(N1670) );
  INVX1 gate210 ( .A(N1202), .Y(N1673) );
  INVX1 gate211 ( .A(N1202), .Y(N1674) );
  INVX1 gate212 ( .A(N1202), .Y(N1675) );
  INVX1 gate213 ( .A(N1202), .Y(N1676) );
  INVX1 gate214 ( .A(N1202), .Y(N1677) );
  INVX1 gate215 ( .A(N1202), .Y(N1678) );
  INVX1 gate216 ( .A(N1202), .Y(N1679) );
  INVX1 gate217 ( .A(N1202), .Y(N1680) );
  NAND2X1 gate218 ( .A(N941), .B(N1467), .Y(N1691) );
  NAND2X1 gate219 ( .A(N938), .B(N1468), .Y(N1692) );
  NAND2X1 gate220 ( .A(N947), .B(N1469), .Y(N1693) );
  NAND2X1 gate221 ( .A(N944), .B(N1470), .Y(N1694) );
  INVX1 gate222 ( .A(N1505), .Y(N1713) );
  AND2X1 gate223 ( .A(N87), .B(N1264), .Y(N1714) );
  NAND2X1 gate224 ( .A(N1509), .B(N1510), .Y(N1715) );
  NAND2X1 gate225 ( .A(N1511), .B(N1512), .Y(N1718) );
  NAND2X1 gate226 ( .A(N1507), .B(N1508), .Y(N1721) );
  AND2X1 gate227 ( .A(N763), .B(N1340), .Y(N1722) );
  NAND2X1 gate228 ( .A(N763), .B(N1340), .Y(N1725) );
  INVX1 gate229 ( .A(N1268), .Y(N1726) );
  NAND2X1 gate230 ( .A(N1493), .B(N1271), .Y(N1727) );
  INVX1 gate231 ( .A(N1493), .Y(N1728) );
  AND2X1 gate232 ( .A(N683), .B(N1268), .Y(N1729) );
  NAND2X1 gate233 ( .A(N1499), .B(N1272), .Y(N1730) );
  INVX1 gate234 ( .A(N1499), .Y(N1731) );
  NAND2X1 gate235 ( .A(N87), .B(N1264), .Y(N1735) );
  INVX1 gate236 ( .A(N1273), .Y(N1736) );
  INVX1 gate237 ( .A(N1276), .Y(N1737) );
  NAND2X1 gate238 ( .A(N1325), .B(N821), .Y(N1738) );
  NAND2X1 gate239 ( .A(N1325), .B(N825), .Y(N1747) );
  NAND3X1 gate240 ( .A(N772), .B(N1279), .C(N798), .Y(N1756) );
  NAND2X1 gate241_1 ( .A(N772), .B(N786), .Y(N1761_1) );
  NAND2X1 gate241_2 ( .A(N798), .B(N1302), .Y(N1761_2) );
  NAND2X1 gate241 ( .A(N1761_1), .B(N1761_2), .Y(N1761) );
  NAND2X1 gate242 ( .A(N1496), .B(N1339), .Y(N1764) );
  INVX1 gate243 ( .A(N1496), .Y(N1765) );
  NAND2X1 gate244 ( .A(N1502), .B(N1344), .Y(N1766) );
  INVX1 gate245 ( .A(N1502), .Y(N1767) );
  INVX1 gate246 ( .A(N1328), .Y(N1768) );
  INVX1 gate247 ( .A(N1334), .Y(N1769) );
  INVX1 gate248 ( .A(N1331), .Y(N1770) );
  AND2X1 gate249 ( .A(N845), .B(N1579), .Y(N1787) );
  AND2X1 gate250 ( .A(N150), .B(N1580), .Y(N1788) );
  AND2X1 gate251 ( .A(N851), .B(N1582), .Y(N1789) );
  AND2X1 gate252 ( .A(N159), .B(N1583), .Y(N1790) );
  AND2X1 gate253 ( .A(N77), .B(N1584), .Y(N1791) );
  AND2X1 gate254 ( .A(N50), .B(N1585), .Y(N1792) );
  AND2X1 gate255 ( .A(N858), .B(N1587), .Y(N1793) );
  AND2X1 gate256 ( .A(N845), .B(N1588), .Y(N1794) );
  AND2X1 gate257 ( .A(N864), .B(N1590), .Y(N1795) );
  AND2X1 gate258 ( .A(N851), .B(N1591), .Y(N1796) );
  AND2X1 gate259 ( .A(N107), .B(N1593), .Y(N1797) );
  AND2X1 gate260 ( .A(N77), .B(N1594), .Y(N1798) );
  AND2X1 gate261 ( .A(N116), .B(N1595), .Y(N1799) );
  AND2X1 gate262 ( .A(N858), .B(N1596), .Y(N1800) );
  AND2X1 gate263 ( .A(N283), .B(N1598), .Y(N1801) );
  AND2X1 gate264 ( .A(N864), .B(N1599), .Y(N1802) );
  AND2X1 gate265 ( .A(N200), .B(N1363), .Y(N1803) );
  AND2X1 gate266 ( .A(N889), .B(N1363), .Y(N1806) );
  AND2X1 gate267 ( .A(N890), .B(N1366), .Y(N1809) );
  AND2X1 gate268 ( .A(N891), .B(N1366), .Y(N1812) );
  NAND2X1 gate269 ( .A(N1298), .B(N1302), .Y(N1815) );
  NAND2X1 gate270 ( .A(N821), .B(N1302), .Y(N1818) );
  NAND3X1 gate271 ( .A(N772), .B(N1279), .C(N1179), .Y(N1821) );
  NAND3X1 gate272 ( .A(N786), .B(N794), .C(N1298), .Y(N1824) );
  NAND2X1 gate273 ( .A(N786), .B(N1298), .Y(N1833) );
  INVX1 gate274 ( .A(N1369), .Y(N1842) );
  INVX1 gate275 ( .A(N1369), .Y(N1843) );
  INVX1 gate276 ( .A(N1369), .Y(N1844) );
  INVX1 gate277 ( .A(N1369), .Y(N1845) );
  INVX1 gate278 ( .A(N1369), .Y(N1846) );
  INVX1 gate279 ( .A(N1369), .Y(N1847) );
  INVX1 gate280 ( .A(N1369), .Y(N1848) );
  INVX1 gate281 ( .A(N1384), .Y(N1849) );
  AND2X1 gate282 ( .A(N1384), .B(N896), .Y(N1850) );
  INVX1 gate283 ( .A(N1384), .Y(N1851) );
  AND2X1 gate284 ( .A(N1384), .B(N896), .Y(N1852) );
  INVX1 gate285 ( .A(N1384), .Y(N1853) );
  AND2X1 gate286 ( .A(N1384), .B(N896), .Y(N1854) );
  INVX1 gate287 ( .A(N1384), .Y(N1855) );
  AND2X1 gate288 ( .A(N1384), .B(N896), .Y(N1856) );
  INVX1 gate289 ( .A(N1384), .Y(N1857) );
  AND2X1 gate290 ( .A(N1384), .B(N896), .Y(N1858) );
  INVX1 gate291 ( .A(N1384), .Y(N1859) );
  AND2X1 gate292 ( .A(N1384), .B(N896), .Y(N1860) );
  INVX1 gate293 ( .A(N1384), .Y(N1861) );
  AND2X1 gate294 ( .A(N1384), .B(N896), .Y(N1862) );
  INVX1 gate295 ( .A(N1384), .Y(N1863) );
  AND2X1 gate296 ( .A(N1384), .B(N896), .Y(N1864) );
  AND2X1 gate297 ( .A(N1202), .B(N1409), .Y(N1869) );
  NOR2X1 gate298 ( .A(N50), .B(N1409), .Y(N1870) );
  INVX1 gate299 ( .A(N1306), .Y(N1873) );
  AND2X1 gate300 ( .A(N1202), .B(N1409), .Y(N1874) );
  NOR2X1 gate301 ( .A(N58), .B(N1409), .Y(N1875) );
  INVX1 gate302 ( .A(N1306), .Y(N1878) );
  AND2X1 gate303 ( .A(N1202), .B(N1409), .Y(N1879) );
  NOR2X1 gate304 ( .A(N68), .B(N1409), .Y(N1880) );
  INVX1 gate305 ( .A(N1306), .Y(N1883) );
  AND2X1 gate306 ( .A(N1202), .B(N1409), .Y(N1884) );
  NOR2X1 gate307 ( .A(N77), .B(N1409), .Y(N1885) );
  INVX1 gate308 ( .A(N1306), .Y(N1888) );
  AND2X1 gate309 ( .A(N1202), .B(N1409), .Y(N1889) );
  NOR2X1 gate310 ( .A(N87), .B(N1409), .Y(N1890) );
  INVX1 gate311 ( .A(N1322), .Y(N1893) );
  AND2X1 gate312 ( .A(N1202), .B(N1409), .Y(N1894) );
  NOR2X1 gate313 ( .A(N97), .B(N1409), .Y(N1895) );
  INVX1 gate314 ( .A(N1315), .Y(N1898) );
  AND2X1 gate315 ( .A(N1202), .B(N1409), .Y(N1899) );
  NOR2X1 gate316 ( .A(N107), .B(N1409), .Y(N1900) );
  INVX1 gate317 ( .A(N1315), .Y(N1903) );
  AND2X1 gate318 ( .A(N1202), .B(N1409), .Y(N1904) );
  NOR2X1 gate319 ( .A(N116), .B(N1409), .Y(N1905) );
  INVX1 gate320 ( .A(N1315), .Y(N1908) );
  AND2X1 gate321 ( .A(N1452), .B(N213), .Y(N1909) );
  NAND2X1 gate322 ( .A(N1452), .B(N213), .Y(N1912) );
  AND2X1 gate323_1 ( .A(N1452), .B(N213), .Y(N1913_1) );
  AND2X1 gate323 ( .A(N343), .B(N1913_1), .Y(N1913) );
  NAND3X1 gate324 ( .A(N1452), .B(N213), .C(N343), .Y(N1917) );
  AND2X1 gate325_1 ( .A(N1452), .B(N213), .Y(N1922_1) );
  AND2X1 gate325 ( .A(N343), .B(N1922_1), .Y(N1922) );
  NAND3X1 gate326 ( .A(N1452), .B(N213), .C(N343), .Y(N1926) );
  BUFX2 gate327 ( .A(N1464), .Y(N1930) );
  NAND2X1 gate328 ( .A(N1691), .B(N1692), .Y(N1933) );
  NAND2X1 gate329 ( .A(N1693), .B(N1694), .Y(N1936) );
  INVX1 gate330 ( .A(N1471), .Y(N1939) );
  NAND2X1 gate331 ( .A(N1471), .B(N1474), .Y(N1940) );
  INVX1 gate332 ( .A(N1475), .Y(N1941) );
  INVX1 gate333 ( .A(N1478), .Y(N1942) );
  INVX1 gate334 ( .A(N1481), .Y(N1943) );
  INVX1 gate335 ( .A(N1484), .Y(N1944) );
  INVX1 gate336 ( .A(N1487), .Y(N1945) );
  INVX1 gate337 ( .A(N1490), .Y(N1946) );
  INVX1 gate338 ( .A(N1714), .Y(N1947) );
  NAND2X1 gate339 ( .A(N953), .B(N1728), .Y(N1960) );
  NAND2X1 gate340 ( .A(N959), .B(N1731), .Y(N1961) );
  AND2X1 gate341 ( .A(N1520), .B(N1276), .Y(N1966) );
  NAND2X1 gate342 ( .A(N956), .B(N1765), .Y(N1981) );
  NAND2X1 gate343 ( .A(N962), .B(N1767), .Y(N1982) );
  AND2X1 gate344 ( .A(N1067), .B(N1768), .Y(N1983) );
  OR2X1 gate345_1 ( .A(N1581), .B(N1787), .Y(N1986_1) );
  OR2X1 gate345 ( .A(N1788), .B(N1986_1), .Y(N1986) );
  OR2X1 gate346_1 ( .A(N1586), .B(N1791), .Y(N1987_1) );
  OR2X1 gate346 ( .A(N1792), .B(N1987_1), .Y(N1987) );
  OR2X1 gate347_1 ( .A(N1589), .B(N1793), .Y(N1988_1) );
  OR2X1 gate347 ( .A(N1794), .B(N1988_1), .Y(N1988) );
  OR2X1 gate348_1 ( .A(N1592), .B(N1795), .Y(N1989_1) );
  OR2X1 gate348 ( .A(N1796), .B(N1989_1), .Y(N1989) );
  OR2X1 gate349_1 ( .A(N1597), .B(N1799), .Y(N1990_1) );
  OR2X1 gate349 ( .A(N1800), .B(N1990_1), .Y(N1990) );
  OR2X1 gate350_1 ( .A(N1600), .B(N1801), .Y(N1991_1) );
  OR2X1 gate350 ( .A(N1802), .B(N1991_1), .Y(N1991) );
  AND2X1 gate351 ( .A(N77), .B(N1849), .Y(N2022) );
  AND2X1 gate352 ( .A(N223), .B(N1850), .Y(N2023) );
  AND2X1 gate353 ( .A(N87), .B(N1851), .Y(N2024) );
  AND2X1 gate354 ( .A(N226), .B(N1852), .Y(N2025) );
  AND2X1 gate355 ( .A(N97), .B(N1853), .Y(N2026) );
  AND2X1 gate356 ( .A(N232), .B(N1854), .Y(N2027) );
  AND2X1 gate357 ( .A(N107), .B(N1855), .Y(N2028) );
  AND2X1 gate358 ( .A(N238), .B(N1856), .Y(N2029) );
  AND2X1 gate359 ( .A(N116), .B(N1857), .Y(N2030) );
  AND2X1 gate360 ( .A(N244), .B(N1858), .Y(N2031) );
  AND2X1 gate361 ( .A(N283), .B(N1859), .Y(N2032) );
  AND2X1 gate362 ( .A(N250), .B(N1860), .Y(N2033) );
  AND2X1 gate363 ( .A(N294), .B(N1861), .Y(N2034) );
  AND2X1 gate364 ( .A(N257), .B(N1862), .Y(N2035) );
  AND2X1 gate365 ( .A(N303), .B(N1863), .Y(N2036) );
  AND2X1 gate366 ( .A(N264), .B(N1864), .Y(N2037) );
  BUFX2 gate367 ( .A(N1667), .Y(N2038) );
  INVX1 gate368 ( .A(N1667), .Y(N2043) );
  BUFX2 gate369 ( .A(N1670), .Y(N2052) );
  INVX1 gate370 ( .A(N1670), .Y(N2057) );
  AND2X1 gate371_1 ( .A(N50), .B(N1197), .Y(N2068_1) );
  AND2X1 gate371 ( .A(N1869), .B(N2068_1), .Y(N2068) );
  AND2X1 gate372_1 ( .A(N58), .B(N1197), .Y(N2073_1) );
  AND2X1 gate372 ( .A(N1874), .B(N2073_1), .Y(N2073) );
  AND2X1 gate373_1 ( .A(N68), .B(N1197), .Y(N2078_1) );
  AND2X1 gate373 ( .A(N1879), .B(N2078_1), .Y(N2078) );
  AND2X1 gate374_1 ( .A(N77), .B(N1197), .Y(N2083_1) );
  AND2X1 gate374 ( .A(N1884), .B(N2083_1), .Y(N2083) );
  AND2X1 gate375_1 ( .A(N87), .B(N1219), .Y(N2088_1) );
  AND2X1 gate375 ( .A(N1889), .B(N2088_1), .Y(N2088) );
  AND2X1 gate376_1 ( .A(N97), .B(N1219), .Y(N2093_1) );
  AND2X1 gate376 ( .A(N1894), .B(N2093_1), .Y(N2093) );
  AND2X1 gate377_1 ( .A(N107), .B(N1219), .Y(N2098_1) );
  AND2X1 gate377 ( .A(N1899), .B(N2098_1), .Y(N2098) );
  AND2X1 gate378_1 ( .A(N116), .B(N1219), .Y(N2103_1) );
  AND2X1 gate378 ( .A(N1904), .B(N2103_1), .Y(N2103) );
  INVX1 gate379 ( .A(N1562), .Y(N2121) );
  INVX1 gate380 ( .A(N1562), .Y(N2122) );
  INVX1 gate381 ( .A(N1562), .Y(N2123) );
  INVX1 gate382 ( .A(N1562), .Y(N2124) );
  INVX1 gate383 ( .A(N1562), .Y(N2125) );
  INVX1 gate384 ( .A(N1562), .Y(N2126) );
  INVX1 gate385 ( .A(N1562), .Y(N2127) );
  INVX1 gate386 ( .A(N1562), .Y(N2128) );
  NAND2X1 gate387 ( .A(N950), .B(N1939), .Y(N2133) );
  NAND2X1 gate388 ( .A(N1478), .B(N1941), .Y(N2134) );
  NAND2X1 gate389 ( .A(N1475), .B(N1942), .Y(N2135) );
  NAND2X1 gate390 ( .A(N1484), .B(N1943), .Y(N2136) );
  NAND2X1 gate391 ( .A(N1481), .B(N1944), .Y(N2137) );
  NAND2X1 gate392 ( .A(N1490), .B(N1945), .Y(N2138) );
  NAND2X1 gate393 ( .A(N1487), .B(N1946), .Y(N2139) );
  INVX1 gate394 ( .A(N1933), .Y(N2141) );
  INVX1 gate395 ( .A(N1936), .Y(N2142) );
  INVX1 gate396 ( .A(N1738), .Y(N2143) );
  AND2X1 gate397 ( .A(N1738), .B(N1747), .Y(N2144) );
  INVX1 gate398 ( .A(N1747), .Y(N2145) );
  NAND2X1 gate399 ( .A(N1727), .B(N1960), .Y(N2146) );
  NAND2X1 gate400 ( .A(N1730), .B(N1961), .Y(N2147) );
  AND2X1 gate401_1 ( .A(N1722), .B(N1267), .Y(N2148_1) );
  AND2X1 gate401_2 ( .A(N665), .B(N58), .Y(N2148_2) );
  AND2X1 gate401 ( .A(N2148_1), .B(N2148_2), .Y(N2148) );
  INVX1 gate402 ( .A(N1738), .Y(N2149) );
  AND2X1 gate403 ( .A(N1738), .B(N1747), .Y(N2150) );
  INVX1 gate404 ( .A(N1747), .Y(N2151) );
  INVX1 gate405 ( .A(N1738), .Y(N2152) );
  INVX1 gate406 ( .A(N1747), .Y(N2153) );
  AND2X1 gate407 ( .A(N1738), .B(N1747), .Y(N2154) );
  INVX1 gate408 ( .A(N1738), .Y(N2155) );
  INVX1 gate409 ( .A(N1747), .Y(N2156) );
  AND2X1 gate410 ( .A(N1738), .B(N1747), .Y(N2157) );
  BUFX2 gate411 ( .A(N1761), .Y(N2158) );
  BUFX2 gate412 ( .A(N1761), .Y(N2175) );
  NAND2X1 gate413 ( .A(N1764), .B(N1981), .Y(N2178) );
  NAND2X1 gate414 ( .A(N1766), .B(N1982), .Y(N2179) );
  INVX1 gate415 ( .A(N1756), .Y(N2180) );
  AND2X1 gate416 ( .A(N1756), .B(N1328), .Y(N2181) );
  INVX1 gate417 ( .A(N1756), .Y(N2183) );
  AND2X1 gate418 ( .A(N1331), .B(N1756), .Y(N2184) );
  NAND2X1 gate419 ( .A(N1358), .B(N1812), .Y(N2185) );
  NAND2X1 gate420 ( .A(N1358), .B(N1809), .Y(N2188) );
  NAND2X1 gate421 ( .A(N1353), .B(N1812), .Y(N2191) );
  NAND2X1 gate422 ( .A(N1353), .B(N1809), .Y(N2194) );
  NAND2X1 gate423 ( .A(N1358), .B(N1806), .Y(N2197) );
  NAND2X1 gate424 ( .A(N1358), .B(N1803), .Y(N2200) );
  NAND2X1 gate425 ( .A(N1353), .B(N1806), .Y(N2203) );
  NAND2X1 gate426 ( .A(N1353), .B(N1803), .Y(N2206) );
  INVX1 gate427 ( .A(N1815), .Y(N2209) );
  INVX1 gate428 ( .A(N1818), .Y(N2210) );
  AND2X1 gate429 ( .A(N1815), .B(N1818), .Y(N2211) );
  BUFX2 gate430 ( .A(N1821), .Y(N2212) );
  BUFX2 gate431 ( .A(N1821), .Y(N2221) );
  INVX1 gate432 ( .A(N1833), .Y(N2230) );
  INVX1 gate433 ( .A(N1833), .Y(N2231) );
  INVX1 gate434 ( .A(N1833), .Y(N2232) );
  INVX1 gate435 ( .A(N1833), .Y(N2233) );
  INVX1 gate436 ( .A(N1824), .Y(N2234) );
  INVX1 gate437 ( .A(N1824), .Y(N2235) );
  INVX1 gate438 ( .A(N1824), .Y(N2236) );
  INVX1 gate439 ( .A(N1824), .Y(N2237) );
  OR2X1 gate440_1 ( .A(N2022), .B(N1643), .Y(N2238_1) );
  OR2X1 gate440 ( .A(N2023), .B(N2238_1), .Y(N2238) );
  OR2X1 gate441_1 ( .A(N2024), .B(N1644), .Y(N2239_1) );
  OR2X1 gate441 ( .A(N2025), .B(N2239_1), .Y(N2239) );
  OR2X1 gate442_1 ( .A(N2026), .B(N1645), .Y(N2240_1) );
  OR2X1 gate442 ( .A(N2027), .B(N2240_1), .Y(N2240) );
  OR2X1 gate443_1 ( .A(N2028), .B(N1646), .Y(N2241_1) );
  OR2X1 gate443 ( .A(N2029), .B(N2241_1), .Y(N2241) );
  OR2X1 gate444_1 ( .A(N2030), .B(N1647), .Y(N2242_1) );
  OR2X1 gate444 ( .A(N2031), .B(N2242_1), .Y(N2242) );
  OR2X1 gate445_1 ( .A(N2032), .B(N1648), .Y(N2243_1) );
  OR2X1 gate445 ( .A(N2033), .B(N2243_1), .Y(N2243) );
  OR2X1 gate446_1 ( .A(N2034), .B(N1649), .Y(N2244_1) );
  OR2X1 gate446 ( .A(N2035), .B(N2244_1), .Y(N2244) );
  OR2X1 gate447_1 ( .A(N2036), .B(N1650), .Y(N2245_1) );
  OR2X1 gate447 ( .A(N2037), .B(N2245_1), .Y(N2245) );
  AND2X1 gate448 ( .A(N1986), .B(N1673), .Y(N2270) );
  AND2X1 gate449 ( .A(N1987), .B(N1675), .Y(N2277) );
  AND2X1 gate450 ( .A(N1988), .B(N1676), .Y(N2282) );
  AND2X1 gate451 ( .A(N1989), .B(N1677), .Y(N2287) );
  AND2X1 gate452 ( .A(N1990), .B(N1679), .Y(N2294) );
  AND2X1 gate453 ( .A(N1991), .B(N1680), .Y(N2299) );
  BUFX2 gate454 ( .A(N1917), .Y(N2304) );
  AND2X1 gate455 ( .A(N1930), .B(N350), .Y(N2307) );
  NAND2X1 gate456 ( .A(N1930), .B(N350), .Y(N2310) );
  BUFX2 gate457 ( .A(N1715), .Y(N2313) );
  BUFX2 gate458 ( .A(N1718), .Y(N2316) );
  BUFX2 gate459 ( .A(N1715), .Y(N2319) );
  BUFX2 gate460 ( .A(N1718), .Y(N2322) );
  NAND2X1 gate461 ( .A(N1940), .B(N2133), .Y(N2325) );
  NAND2X1 gate462 ( .A(N2134), .B(N2135), .Y(N2328) );
  NAND2X1 gate463 ( .A(N2136), .B(N2137), .Y(N2331) );
  NAND2X1 gate464 ( .A(N2138), .B(N2139), .Y(N2334) );
  NAND2X1 gate465 ( .A(N1936), .B(N2141), .Y(N2341) );
  NAND2X1 gate466 ( .A(N1933), .B(N2142), .Y(N2342) );
  AND2X1 gate467 ( .A(N724), .B(N2144), .Y(N2347) );
  AND2X1 gate468_1 ( .A(N2146), .B(N699), .Y(N2348_1) );
  AND2X1 gate468 ( .A(N1726), .B(N2348_1), .Y(N2348) );
  AND2X1 gate469 ( .A(N753), .B(N2147), .Y(N2349) );
  AND2X1 gate470 ( .A(N2148), .B(N1273), .Y(N2350) );
  AND2X1 gate471 ( .A(N736), .B(N2150), .Y(N2351) );
  AND2X1 gate472 ( .A(N1735), .B(N2153), .Y(N2352) );
  AND2X1 gate473 ( .A(N763), .B(N2154), .Y(N2353) );
  AND2X1 gate474 ( .A(N1725), .B(N2156), .Y(N2354) );
  AND2X1 gate475 ( .A(N749), .B(N2157), .Y(N2355) );
  INVX1 gate476 ( .A(N2178), .Y(N2374) );
  INVX1 gate477 ( .A(N2179), .Y(N2375) );
  AND2X1 gate478 ( .A(N1520), .B(N2180), .Y(N2376) );
  AND2X1 gate479 ( .A(N1721), .B(N2181), .Y(N2379) );
  AND2X1 gate480 ( .A(N665), .B(N2211), .Y(N2398) );
  AND2X1 gate481_1 ( .A(N2057), .B(N226), .Y(N2417_1) );
  AND2X1 gate481 ( .A(N1873), .B(N2417_1), .Y(N2417) );
  AND2X1 gate482_1 ( .A(N2057), .B(N274), .Y(N2418_1) );
  AND2X1 gate482 ( .A(N1306), .B(N2418_1), .Y(N2418) );
  AND2X1 gate483 ( .A(N2052), .B(N2238), .Y(N2419) );
  AND2X1 gate484_1 ( .A(N2057), .B(N232), .Y(N2420_1) );
  AND2X1 gate484 ( .A(N1878), .B(N2420_1), .Y(N2420) );
  AND2X1 gate485_1 ( .A(N2057), .B(N274), .Y(N2421_1) );
  AND2X1 gate485 ( .A(N1306), .B(N2421_1), .Y(N2421) );
  AND2X1 gate486 ( .A(N2052), .B(N2239), .Y(N2422) );
  AND2X1 gate487_1 ( .A(N2057), .B(N238), .Y(N2425_1) );
  AND2X1 gate487 ( .A(N1883), .B(N2425_1), .Y(N2425) );
  AND2X1 gate488_1 ( .A(N2057), .B(N274), .Y(N2426_1) );
  AND2X1 gate488 ( .A(N1306), .B(N2426_1), .Y(N2426) );
  AND2X1 gate489 ( .A(N2052), .B(N2240), .Y(N2427) );
  AND2X1 gate490_1 ( .A(N2057), .B(N244), .Y(N2430_1) );
  AND2X1 gate490 ( .A(N1888), .B(N2430_1), .Y(N2430) );
  AND2X1 gate491_1 ( .A(N2057), .B(N274), .Y(N2431_1) );
  AND2X1 gate491 ( .A(N1306), .B(N2431_1), .Y(N2431) );
  AND2X1 gate492 ( .A(N2052), .B(N2241), .Y(N2432) );
  AND2X1 gate493_1 ( .A(N2043), .B(N250), .Y(N2435_1) );
  AND2X1 gate493 ( .A(N1893), .B(N2435_1), .Y(N2435) );
  AND2X1 gate494_1 ( .A(N2043), .B(N274), .Y(N2436_1) );
  AND2X1 gate494 ( .A(N1322), .B(N2436_1), .Y(N2436) );
  AND2X1 gate495 ( .A(N2038), .B(N2242), .Y(N2437) );
  AND2X1 gate496_1 ( .A(N2043), .B(N257), .Y(N2438_1) );
  AND2X1 gate496 ( .A(N1898), .B(N2438_1), .Y(N2438) );
  AND2X1 gate497_1 ( .A(N2043), .B(N274), .Y(N2439_1) );
  AND2X1 gate497 ( .A(N1315), .B(N2439_1), .Y(N2439) );
  AND2X1 gate498 ( .A(N2038), .B(N2243), .Y(N2440) );
  AND2X1 gate499_1 ( .A(N2043), .B(N264), .Y(N2443_1) );
  AND2X1 gate499 ( .A(N1903), .B(N2443_1), .Y(N2443) );
  AND2X1 gate500_1 ( .A(N2043), .B(N274), .Y(N2444_1) );
  AND2X1 gate500 ( .A(N1315), .B(N2444_1), .Y(N2444) );
  AND2X1 gate501 ( .A(N2038), .B(N2244), .Y(N2445) );
  AND2X1 gate502_1 ( .A(N2043), .B(N270), .Y(N2448_1) );
  AND2X1 gate502 ( .A(N1908), .B(N2448_1), .Y(N2448) );
  AND2X1 gate503_1 ( .A(N2043), .B(N274), .Y(N2449_1) );
  AND2X1 gate503 ( .A(N1315), .B(N2449_1), .Y(N2449) );
  AND2X1 gate504 ( .A(N2038), .B(N2245), .Y(N2450) );
  INVX1 gate505 ( .A(N2313), .Y(N2467) );
  INVX1 gate506 ( .A(N2316), .Y(N2468) );
  INVX1 gate507 ( .A(N2319), .Y(N2469) );
  INVX1 gate508 ( .A(N2322), .Y(N2470) );
  NAND2X1 gate509 ( .A(N2341), .B(N2342), .Y(N2471) );
  INVX1 gate510 ( .A(N2325), .Y(N2474) );
  INVX1 gate511 ( .A(N2328), .Y(N2475) );
  INVX1 gate512 ( .A(N2331), .Y(N2476) );
  INVX1 gate513 ( .A(N2334), .Y(N2477) );
  OR2X1 gate514 ( .A(N2348), .B(N1729), .Y(N2478) );
  INVX1 gate515 ( .A(N2175), .Y(N2481) );
  AND2X1 gate516 ( .A(N2175), .B(N1334), .Y(N2482) );
  AND2X1 gate517 ( .A(N2349), .B(N2183), .Y(N2483) );
  AND2X1 gate518 ( .A(N2374), .B(N1346), .Y(N2486) );
  AND2X1 gate519 ( .A(N2375), .B(N1350), .Y(N2487) );
  BUFX2 gate520 ( .A(N2185), .Y(N2488) );
  BUFX2 gate521 ( .A(N2188), .Y(N2497) );
  BUFX2 gate522 ( .A(N2191), .Y(N2506) );
  BUFX2 gate523 ( .A(N2194), .Y(N2515) );
  BUFX2 gate524 ( .A(N2197), .Y(N2524) );
  BUFX2 gate525 ( .A(N2200), .Y(N2533) );
  BUFX2 gate526 ( .A(N2203), .Y(N2542) );
  BUFX2 gate527 ( .A(N2206), .Y(N2551) );
  BUFX2 gate528 ( .A(N2185), .Y(N2560) );
  BUFX2 gate529 ( .A(N2188), .Y(N2569) );
  BUFX2 gate530 ( .A(N2191), .Y(N2578) );
  BUFX2 gate531 ( .A(N2194), .Y(N2587) );
  BUFX2 gate532 ( .A(N2197), .Y(N2596) );
  BUFX2 gate533 ( .A(N2200), .Y(N2605) );
  BUFX2 gate534 ( .A(N2203), .Y(N2614) );
  BUFX2 gate535 ( .A(N2206), .Y(N2623) );
  INVX1 gate536 ( .A(N2212), .Y(N2632) );
  AND2X1 gate537 ( .A(N2212), .B(N1833), .Y(N2633) );
  INVX1 gate538 ( .A(N2212), .Y(N2634) );
  AND2X1 gate539 ( .A(N2212), .B(N1833), .Y(N2635) );
  INVX1 gate540 ( .A(N2212), .Y(N2636) );
  AND2X1 gate541 ( .A(N2212), .B(N1833), .Y(N2637) );
  INVX1 gate542 ( .A(N2212), .Y(N2638) );
  AND2X1 gate543 ( .A(N2212), .B(N1833), .Y(N2639) );
  INVX1 gate544 ( .A(N2221), .Y(N2640) );
  AND2X1 gate545 ( .A(N2221), .B(N1824), .Y(N2641) );
  INVX1 gate546 ( .A(N2221), .Y(N2642) );
  AND2X1 gate547 ( .A(N2221), .B(N1824), .Y(N2643) );
  INVX1 gate548 ( .A(N2221), .Y(N2644) );
  AND2X1 gate549 ( .A(N2221), .B(N1824), .Y(N2645) );
  INVX1 gate550 ( .A(N2221), .Y(N2646) );
  AND2X1 gate551 ( .A(N2221), .B(N1824), .Y(N2647) );
  OR2X1 gate552_1 ( .A(N2270), .B(N1870), .Y(N2648_1) );
  OR2X1 gate552 ( .A(N2068), .B(N2648_1), .Y(N2648) );
  NOR3X1 gate553 ( .A(N2270), .B(N1870), .C(N2068), .Y(N2652) );
  OR2X1 gate554_1 ( .A(N2417), .B(N2418), .Y(N2656_1) );
  OR2X1 gate554 ( .A(N2419), .B(N2656_1), .Y(N2656) );
  OR2X1 gate555_1 ( .A(N2420), .B(N2421), .Y(N2659_1) );
  OR2X1 gate555 ( .A(N2422), .B(N2659_1), .Y(N2659) );
  OR2X1 gate556_1 ( .A(N2277), .B(N1880), .Y(N2662_1) );
  OR2X1 gate556 ( .A(N2078), .B(N2662_1), .Y(N2662) );
  NOR3X1 gate557 ( .A(N2277), .B(N1880), .C(N2078), .Y(N2666) );
  OR2X1 gate558_1 ( .A(N2425), .B(N2426), .Y(N2670_1) );
  OR2X1 gate558 ( .A(N2427), .B(N2670_1), .Y(N2670) );
  OR2X1 gate559_1 ( .A(N2282), .B(N1885), .Y(N2673_1) );
  OR2X1 gate559 ( .A(N2083), .B(N2673_1), .Y(N2673) );
  NOR3X1 gate560 ( .A(N2282), .B(N1885), .C(N2083), .Y(N2677) );
  OR2X1 gate561_1 ( .A(N2430), .B(N2431), .Y(N2681_1) );
  OR2X1 gate561 ( .A(N2432), .B(N2681_1), .Y(N2681) );
  OR2X1 gate562_1 ( .A(N2287), .B(N1890), .Y(N2684_1) );
  OR2X1 gate562 ( .A(N2088), .B(N2684_1), .Y(N2684) );
  NOR3X1 gate563 ( .A(N2287), .B(N1890), .C(N2088), .Y(N2688) );
  OR2X1 gate564_1 ( .A(N2435), .B(N2436), .Y(N2692_1) );
  OR2X1 gate564 ( .A(N2437), .B(N2692_1), .Y(N2692) );
  OR2X1 gate565_1 ( .A(N2438), .B(N2439), .Y(N2697_1) );
  OR2X1 gate565 ( .A(N2440), .B(N2697_1), .Y(N2697) );
  OR2X1 gate566_1 ( .A(N2294), .B(N1900), .Y(N2702_1) );
  OR2X1 gate566 ( .A(N2098), .B(N2702_1), .Y(N2702) );
  NOR3X1 gate567 ( .A(N2294), .B(N1900), .C(N2098), .Y(N2706) );
  OR2X1 gate568_1 ( .A(N2443), .B(N2444), .Y(N2710_1) );
  OR2X1 gate568 ( .A(N2445), .B(N2710_1), .Y(N2710) );
  OR2X1 gate569_1 ( .A(N2299), .B(N1905), .Y(N2715_1) );
  OR2X1 gate569 ( .A(N2103), .B(N2715_1), .Y(N2715) );
  NOR3X1 gate570 ( .A(N2299), .B(N1905), .C(N2103), .Y(N2719) );
  OR2X1 gate571_1 ( .A(N2448), .B(N2449), .Y(N2723_1) );
  OR2X1 gate571 ( .A(N2450), .B(N2723_1), .Y(N2723) );
  INVX1 gate572 ( .A(N2304), .Y(N2728) );
  INVX1 gate573 ( .A(N2158), .Y(N2729) );
  AND2X1 gate574 ( .A(N1562), .B(N2158), .Y(N2730) );
  INVX1 gate575 ( .A(N2158), .Y(N2731) );
  AND2X1 gate576 ( .A(N1562), .B(N2158), .Y(N2732) );
  INVX1 gate577 ( .A(N2158), .Y(N2733) );
  AND2X1 gate578 ( .A(N1562), .B(N2158), .Y(N2734) );
  INVX1 gate579 ( .A(N2158), .Y(N2735) );
  AND2X1 gate580 ( .A(N1562), .B(N2158), .Y(N2736) );
  INVX1 gate581 ( .A(N2158), .Y(N2737) );
  AND2X1 gate582 ( .A(N1562), .B(N2158), .Y(N2738) );
  INVX1 gate583 ( .A(N2158), .Y(N2739) );
  AND2X1 gate584 ( .A(N1562), .B(N2158), .Y(N2740) );
  INVX1 gate585 ( .A(N2158), .Y(N2741) );
  AND2X1 gate586 ( .A(N1562), .B(N2158), .Y(N2742) );
  INVX1 gate587 ( .A(N2158), .Y(N2743) );
  AND2X1 gate588 ( .A(N1562), .B(N2158), .Y(N2744) );
  OR2X1 gate589_1 ( .A(N2376), .B(N1983), .Y(N2745_1) );
  OR2X1 gate589 ( .A(N2379), .B(N2745_1), .Y(N2745) );
  NOR3X1 gate590 ( .A(N2376), .B(N1983), .C(N2379), .Y(N2746) );
  NAND2X1 gate591 ( .A(N2316), .B(N2467), .Y(N2748) );
  NAND2X1 gate592 ( .A(N2313), .B(N2468), .Y(N2749) );
  NAND2X1 gate593 ( .A(N2322), .B(N2469), .Y(N2750) );
  NAND2X1 gate594 ( .A(N2319), .B(N2470), .Y(N2751) );
  NAND2X1 gate595 ( .A(N2328), .B(N2474), .Y(N2754) );
  NAND2X1 gate596 ( .A(N2325), .B(N2475), .Y(N2755) );
  NAND2X1 gate597 ( .A(N2334), .B(N2476), .Y(N2756) );
  NAND2X1 gate598 ( .A(N2331), .B(N2477), .Y(N2757) );
  AND2X1 gate599 ( .A(N1520), .B(N2481), .Y(N2758) );
  AND2X1 gate600 ( .A(N1722), .B(N2482), .Y(N2761) );
  AND2X1 gate601 ( .A(N2478), .B(N1770), .Y(N2764) );
  OR2X1 gate602_1 ( .A(N2486), .B(N1789), .Y(N2768_1) );
  OR2X1 gate602 ( .A(N1790), .B(N2768_1), .Y(N2768) );
  OR2X1 gate603_1 ( .A(N2487), .B(N1797), .Y(N2769_1) );
  OR2X1 gate603 ( .A(N1798), .B(N2769_1), .Y(N2769) );
  AND2X1 gate604 ( .A(N665), .B(N2633), .Y(N2898) );
  AND2X1 gate605 ( .A(N679), .B(N2635), .Y(N2899) );
  AND2X1 gate606 ( .A(N686), .B(N2637), .Y(N2900) );
  AND2X1 gate607 ( .A(N702), .B(N2639), .Y(N2901) );
  INVX1 gate608 ( .A(N2746), .Y(N2962) );
  NAND2X1 gate609 ( .A(N2748), .B(N2749), .Y(N2966) );
  NAND2X1 gate610 ( .A(N2750), .B(N2751), .Y(N2967) );
  BUFX2 gate611 ( .A(N2471), .Y(N2970) );
  NAND2X1 gate612 ( .A(N2754), .B(N2755), .Y(N2973) );
  NAND2X1 gate613 ( .A(N2756), .B(N2757), .Y(N2977) );
  AND2X1 gate614 ( .A(N2471), .B(N2143), .Y(N2980) );
  INVX1 gate615 ( .A(N2488), .Y(N2984) );
  INVX1 gate616 ( .A(N2497), .Y(N2985) );
  INVX1 gate617 ( .A(N2506), .Y(N2986) );
  INVX1 gate618 ( .A(N2515), .Y(N2987) );
  INVX1 gate619 ( .A(N2524), .Y(N2988) );
  INVX1 gate620 ( .A(N2533), .Y(N2989) );
  INVX1 gate621 ( .A(N2542), .Y(N2990) );
  INVX1 gate622 ( .A(N2551), .Y(N2991) );
  INVX1 gate623 ( .A(N2488), .Y(N2992) );
  INVX1 gate624 ( .A(N2497), .Y(N2993) );
  INVX1 gate625 ( .A(N2506), .Y(N2994) );
  INVX1 gate626 ( .A(N2515), .Y(N2995) );
  INVX1 gate627 ( .A(N2524), .Y(N2996) );
  INVX1 gate628 ( .A(N2533), .Y(N2997) );
  INVX1 gate629 ( .A(N2542), .Y(N2998) );
  INVX1 gate630 ( .A(N2551), .Y(N2999) );
  INVX1 gate631 ( .A(N2488), .Y(N3000) );
  INVX1 gate632 ( .A(N2497), .Y(N3001) );
  INVX1 gate633 ( .A(N2506), .Y(N3002) );
  INVX1 gate634 ( .A(N2515), .Y(N3003) );
  INVX1 gate635 ( .A(N2524), .Y(N3004) );
  INVX1 gate636 ( .A(N2533), .Y(N3005) );
  INVX1 gate637 ( .A(N2542), .Y(N3006) );
  INVX1 gate638 ( .A(N2551), .Y(N3007) );
  INVX1 gate639 ( .A(N2488), .Y(N3008) );
  INVX1 gate640 ( .A(N2497), .Y(N3009) );
  INVX1 gate641 ( .A(N2506), .Y(N3010) );
  INVX1 gate642 ( .A(N2515), .Y(N3011) );
  INVX1 gate643 ( .A(N2524), .Y(N3012) );
  INVX1 gate644 ( .A(N2533), .Y(N3013) );
  INVX1 gate645 ( .A(N2542), .Y(N3014) );
  INVX1 gate646 ( .A(N2551), .Y(N3015) );
  INVX1 gate647 ( .A(N2488), .Y(N3016) );
  INVX1 gate648 ( .A(N2497), .Y(N3017) );
  INVX1 gate649 ( .A(N2506), .Y(N3018) );
  INVX1 gate650 ( .A(N2515), .Y(N3019) );
  INVX1 gate651 ( .A(N2524), .Y(N3020) );
  INVX1 gate652 ( .A(N2533), .Y(N3021) );
  INVX1 gate653 ( .A(N2542), .Y(N3022) );
  INVX1 gate654 ( .A(N2551), .Y(N3023) );
  INVX1 gate655 ( .A(N2488), .Y(N3024) );
  INVX1 gate656 ( .A(N2497), .Y(N3025) );
  INVX1 gate657 ( .A(N2506), .Y(N3026) );
  INVX1 gate658 ( .A(N2515), .Y(N3027) );
  INVX1 gate659 ( .A(N2524), .Y(N3028) );
  INVX1 gate660 ( .A(N2533), .Y(N3029) );
  INVX1 gate661 ( .A(N2542), .Y(N3030) );
  INVX1 gate662 ( .A(N2551), .Y(N3031) );
  INVX1 gate663 ( .A(N2488), .Y(N3032) );
  INVX1 gate664 ( .A(N2497), .Y(N3033) );
  INVX1 gate665 ( .A(N2506), .Y(N3034) );
  INVX1 gate666 ( .A(N2515), .Y(N3035) );
  INVX1 gate667 ( .A(N2524), .Y(N3036) );
  INVX1 gate668 ( .A(N2533), .Y(N3037) );
  INVX1 gate669 ( .A(N2542), .Y(N3038) );
  INVX1 gate670 ( .A(N2551), .Y(N3039) );
  INVX1 gate671 ( .A(N2488), .Y(N3040) );
  INVX1 gate672 ( .A(N2497), .Y(N3041) );
  INVX1 gate673 ( .A(N2506), .Y(N3042) );
  INVX1 gate674 ( .A(N2515), .Y(N3043) );
  INVX1 gate675 ( .A(N2524), .Y(N3044) );
  INVX1 gate676 ( .A(N2533), .Y(N3045) );
  INVX1 gate677 ( .A(N2542), .Y(N3046) );
  INVX1 gate678 ( .A(N2551), .Y(N3047) );
  INVX1 gate679 ( .A(N2560), .Y(N3048) );
  INVX1 gate680 ( .A(N2569), .Y(N3049) );
  INVX1 gate681 ( .A(N2578), .Y(N3050) );
  INVX1 gate682 ( .A(N2587), .Y(N3051) );
  INVX1 gate683 ( .A(N2596), .Y(N3052) );
  INVX1 gate684 ( .A(N2605), .Y(N3053) );
  INVX1 gate685 ( .A(N2614), .Y(N3054) );
  INVX1 gate686 ( .A(N2623), .Y(N3055) );
  INVX1 gate687 ( .A(N2560), .Y(N3056) );
  INVX1 gate688 ( .A(N2569), .Y(N3057) );
  INVX1 gate689 ( .A(N2578), .Y(N3058) );
  INVX1 gate690 ( .A(N2587), .Y(N3059) );
  INVX1 gate691 ( .A(N2596), .Y(N3060) );
  INVX1 gate692 ( .A(N2605), .Y(N3061) );
  INVX1 gate693 ( .A(N2614), .Y(N3062) );
  INVX1 gate694 ( .A(N2623), .Y(N3063) );
  INVX1 gate695 ( .A(N2560), .Y(N3064) );
  INVX1 gate696 ( .A(N2569), .Y(N3065) );
  INVX1 gate697 ( .A(N2578), .Y(N3066) );
  INVX1 gate698 ( .A(N2587), .Y(N3067) );
  INVX1 gate699 ( .A(N2596), .Y(N3068) );
  INVX1 gate700 ( .A(N2605), .Y(N3069) );
  INVX1 gate701 ( .A(N2614), .Y(N3070) );
  INVX1 gate702 ( .A(N2623), .Y(N3071) );
  INVX1 gate703 ( .A(N2560), .Y(N3072) );
  INVX1 gate704 ( .A(N2569), .Y(N3073) );
  INVX1 gate705 ( .A(N2578), .Y(N3074) );
  INVX1 gate706 ( .A(N2587), .Y(N3075) );
  INVX1 gate707 ( .A(N2596), .Y(N3076) );
  INVX1 gate708 ( .A(N2605), .Y(N3077) );
  INVX1 gate709 ( .A(N2614), .Y(N3078) );
  INVX1 gate710 ( .A(N2623), .Y(N3079) );
  INVX1 gate711 ( .A(N2560), .Y(N3080) );
  INVX1 gate712 ( .A(N2569), .Y(N3081) );
  INVX1 gate713 ( .A(N2578), .Y(N3082) );
  INVX1 gate714 ( .A(N2587), .Y(N3083) );
  INVX1 gate715 ( .A(N2596), .Y(N3084) );
  INVX1 gate716 ( .A(N2605), .Y(N3085) );
  INVX1 gate717 ( .A(N2614), .Y(N3086) );
  INVX1 gate718 ( .A(N2623), .Y(N3087) );
  INVX1 gate719 ( .A(N2560), .Y(N3088) );
  INVX1 gate720 ( .A(N2569), .Y(N3089) );
  INVX1 gate721 ( .A(N2578), .Y(N3090) );
  INVX1 gate722 ( .A(N2587), .Y(N3091) );
  INVX1 gate723 ( .A(N2596), .Y(N3092) );
  INVX1 gate724 ( .A(N2605), .Y(N3093) );
  INVX1 gate725 ( .A(N2614), .Y(N3094) );
  INVX1 gate726 ( .A(N2623), .Y(N3095) );
  INVX1 gate727 ( .A(N2560), .Y(N3096) );
  INVX1 gate728 ( .A(N2569), .Y(N3097) );
  INVX1 gate729 ( .A(N2578), .Y(N3098) );
  INVX1 gate730 ( .A(N2587), .Y(N3099) );
  INVX1 gate731 ( .A(N2596), .Y(N3100) );
  INVX1 gate732 ( .A(N2605), .Y(N3101) );
  INVX1 gate733 ( .A(N2614), .Y(N3102) );
  INVX1 gate734 ( .A(N2623), .Y(N3103) );
  INVX1 gate735 ( .A(N2560), .Y(N3104) );
  INVX1 gate736 ( .A(N2569), .Y(N3105) );
  INVX1 gate737 ( .A(N2578), .Y(N3106) );
  INVX1 gate738 ( .A(N2587), .Y(N3107) );
  INVX1 gate739 ( .A(N2596), .Y(N3108) );
  INVX1 gate740 ( .A(N2605), .Y(N3109) );
  INVX1 gate741 ( .A(N2614), .Y(N3110) );
  INVX1 gate742 ( .A(N2623), .Y(N3111) );
  BUFX2 gate743 ( .A(N2656), .Y(N3112) );
  INVX1 gate744 ( .A(N2656), .Y(N3115) );
  INVX1 gate745 ( .A(N2652), .Y(N3118) );
  AND2X1 gate746 ( .A(N2768), .B(N1674), .Y(N3119) );
  BUFX2 gate747 ( .A(N2659), .Y(N3122) );
  INVX1 gate748 ( .A(N2659), .Y(N3125) );
  BUFX2 gate749 ( .A(N2670), .Y(N3128) );
  INVX1 gate750 ( .A(N2670), .Y(N3131) );
  INVX1 gate751 ( .A(N2666), .Y(N3134) );
  BUFX2 gate752 ( .A(N2681), .Y(N3135) );
  INVX1 gate753 ( .A(N2681), .Y(N3138) );
  INVX1 gate754 ( .A(N2677), .Y(N3141) );
  BUFX2 gate755 ( .A(N2692), .Y(N3142) );
  INVX1 gate756 ( .A(N2692), .Y(N3145) );
  INVX1 gate757 ( .A(N2688), .Y(N3148) );
  AND2X1 gate758 ( .A(N2769), .B(N1678), .Y(N3149) );
  BUFX2 gate759 ( .A(N2697), .Y(N3152) );
  INVX1 gate760 ( .A(N2697), .Y(N3155) );
  BUFX2 gate761 ( .A(N2710), .Y(N3158) );
  INVX1 gate762 ( .A(N2710), .Y(N3161) );
  INVX1 gate763 ( .A(N2706), .Y(N3164) );
  BUFX2 gate764 ( .A(N2723), .Y(N3165) );
  INVX1 gate765 ( .A(N2723), .Y(N3168) );
  INVX1 gate766 ( .A(N2719), .Y(N3171) );
  AND2X1 gate767 ( .A(N1909), .B(N2648), .Y(N3172) );
  AND2X1 gate768 ( .A(N1913), .B(N2662), .Y(N3175) );
  AND2X1 gate769 ( .A(N1913), .B(N2673), .Y(N3178) );
  AND2X1 gate770 ( .A(N1913), .B(N2684), .Y(N3181) );
  AND2X1 gate771 ( .A(N1922), .B(N2702), .Y(N3184) );
  AND2X1 gate772 ( .A(N1922), .B(N2715), .Y(N3187) );
  INVX1 gate773 ( .A(N2692), .Y(N3190) );
  INVX1 gate774 ( .A(N2697), .Y(N3191) );
  INVX1 gate775 ( .A(N2710), .Y(N3192) );
  INVX1 gate776 ( .A(N2723), .Y(N3193) );
  AND2X1 gate777_1 ( .A(N2692), .B(N2697), .Y(N3194_1) );
  AND2X1 gate777_2 ( .A(N2710), .B(N2723), .Y(N3194_2) );
  AND2X1 gate777_3 ( .A(N1459), .B(N3194_1), .Y(N3194_3) );
  AND2X1 gate777 ( .A(N3194_2), .B(N3194_3), .Y(N3194) );
  NAND2X1 gate778 ( .A(N2745), .B(N2962), .Y(N3195) );
  INVX1 gate779 ( .A(N2966), .Y(N3196) );
  OR2X1 gate780_1 ( .A(N2980), .B(N2145), .Y(N3206_1) );
  OR2X1 gate780 ( .A(N2347), .B(N3206_1), .Y(N3206) );
  AND2X1 gate781 ( .A(N124), .B(N2984), .Y(N3207) );
  AND2X1 gate782 ( .A(N159), .B(N2985), .Y(N3208) );
  AND2X1 gate783 ( .A(N150), .B(N2986), .Y(N3209) );
  AND2X1 gate784 ( .A(N143), .B(N2987), .Y(N3210) );
  AND2X1 gate785 ( .A(N137), .B(N2988), .Y(N3211) );
  AND2X1 gate786 ( .A(N132), .B(N2989), .Y(N3212) );
  AND2X1 gate787 ( .A(N128), .B(N2990), .Y(N3213) );
  AND2X1 gate788 ( .A(N125), .B(N2991), .Y(N3214) );
  AND2X1 gate789 ( .A(N125), .B(N2992), .Y(N3215) );
  AND2X1 gate790 ( .A(N655), .B(N2993), .Y(N3216) );
  AND2X1 gate791 ( .A(N159), .B(N2994), .Y(N3217) );
  AND2X1 gate792 ( .A(N150), .B(N2995), .Y(N3218) );
  AND2X1 gate793 ( .A(N143), .B(N2996), .Y(N3219) );
  AND2X1 gate794 ( .A(N137), .B(N2997), .Y(N3220) );
  AND2X1 gate795 ( .A(N132), .B(N2998), .Y(N3221) );
  AND2X1 gate796 ( .A(N128), .B(N2999), .Y(N3222) );
  AND2X1 gate797 ( .A(N128), .B(N3000), .Y(N3223) );
  AND2X1 gate798 ( .A(N670), .B(N3001), .Y(N3224) );
  AND2X1 gate799 ( .A(N655), .B(N3002), .Y(N3225) );
  AND2X1 gate800 ( .A(N159), .B(N3003), .Y(N3226) );
  AND2X1 gate801 ( .A(N150), .B(N3004), .Y(N3227) );
  AND2X1 gate802 ( .A(N143), .B(N3005), .Y(N3228) );
  AND2X1 gate803 ( .A(N137), .B(N3006), .Y(N3229) );
  AND2X1 gate804 ( .A(N132), .B(N3007), .Y(N3230) );
  AND2X1 gate805 ( .A(N132), .B(N3008), .Y(N3231) );
  AND2X1 gate806 ( .A(N690), .B(N3009), .Y(N3232) );
  AND2X1 gate807 ( .A(N670), .B(N3010), .Y(N3233) );
  AND2X1 gate808 ( .A(N655), .B(N3011), .Y(N3234) );
  AND2X1 gate809 ( .A(N159), .B(N3012), .Y(N3235) );
  AND2X1 gate810 ( .A(N150), .B(N3013), .Y(N3236) );
  AND2X1 gate811 ( .A(N143), .B(N3014), .Y(N3237) );
  AND2X1 gate812 ( .A(N137), .B(N3015), .Y(N3238) );
  AND2X1 gate813 ( .A(N137), .B(N3016), .Y(N3239) );
  AND2X1 gate814 ( .A(N706), .B(N3017), .Y(N3240) );
  AND2X1 gate815 ( .A(N690), .B(N3018), .Y(N3241) );
  AND2X1 gate816 ( .A(N670), .B(N3019), .Y(N3242) );
  AND2X1 gate817 ( .A(N655), .B(N3020), .Y(N3243) );
  AND2X1 gate818 ( .A(N159), .B(N3021), .Y(N3244) );
  AND2X1 gate819 ( .A(N150), .B(N3022), .Y(N3245) );
  AND2X1 gate820 ( .A(N143), .B(N3023), .Y(N3246) );
  AND2X1 gate821 ( .A(N143), .B(N3024), .Y(N3247) );
  AND2X1 gate822 ( .A(N715), .B(N3025), .Y(N3248) );
  AND2X1 gate823 ( .A(N706), .B(N3026), .Y(N3249) );
  AND2X1 gate824 ( .A(N690), .B(N3027), .Y(N3250) );
  AND2X1 gate825 ( .A(N670), .B(N3028), .Y(N3251) );
  AND2X1 gate826 ( .A(N655), .B(N3029), .Y(N3252) );
  AND2X1 gate827 ( .A(N159), .B(N3030), .Y(N3253) );
  AND2X1 gate828 ( .A(N150), .B(N3031), .Y(N3254) );
  AND2X1 gate829 ( .A(N150), .B(N3032), .Y(N3255) );
  AND2X1 gate830 ( .A(N727), .B(N3033), .Y(N3256) );
  AND2X1 gate831 ( .A(N715), .B(N3034), .Y(N3257) );
  AND2X1 gate832 ( .A(N706), .B(N3035), .Y(N3258) );
  AND2X1 gate833 ( .A(N690), .B(N3036), .Y(N3259) );
  AND2X1 gate834 ( .A(N670), .B(N3037), .Y(N3260) );
  AND2X1 gate835 ( .A(N655), .B(N3038), .Y(N3261) );
  AND2X1 gate836 ( .A(N159), .B(N3039), .Y(N3262) );
  AND2X1 gate837 ( .A(N159), .B(N3040), .Y(N3263) );
  AND2X1 gate838 ( .A(N740), .B(N3041), .Y(N3264) );
  AND2X1 gate839 ( .A(N727), .B(N3042), .Y(N3265) );
  AND2X1 gate840 ( .A(N715), .B(N3043), .Y(N3266) );
  AND2X1 gate841 ( .A(N706), .B(N3044), .Y(N3267) );
  AND2X1 gate842 ( .A(N690), .B(N3045), .Y(N3268) );
  AND2X1 gate843 ( .A(N670), .B(N3046), .Y(N3269) );
  AND2X1 gate844 ( .A(N655), .B(N3047), .Y(N3270) );
  AND2X1 gate845 ( .A(N283), .B(N3048), .Y(N3271) );
  AND2X1 gate846 ( .A(N670), .B(N3049), .Y(N3272) );
  AND2X1 gate847 ( .A(N690), .B(N3050), .Y(N3273) );
  AND2X1 gate848 ( .A(N706), .B(N3051), .Y(N3274) );
  AND2X1 gate849 ( .A(N715), .B(N3052), .Y(N3275) );
  AND2X1 gate850 ( .A(N727), .B(N3053), .Y(N3276) );
  AND2X1 gate851 ( .A(N740), .B(N3054), .Y(N3277) );
  AND2X1 gate852 ( .A(N753), .B(N3055), .Y(N3278) );
  AND2X1 gate853 ( .A(N294), .B(N3056), .Y(N3279) );
  AND2X1 gate854 ( .A(N690), .B(N3057), .Y(N3280) );
  AND2X1 gate855 ( .A(N706), .B(N3058), .Y(N3281) );
  AND2X1 gate856 ( .A(N715), .B(N3059), .Y(N3282) );
  AND2X1 gate857 ( .A(N727), .B(N3060), .Y(N3283) );
  AND2X1 gate858 ( .A(N740), .B(N3061), .Y(N3284) );
  AND2X1 gate859 ( .A(N753), .B(N3062), .Y(N3285) );
  AND2X1 gate860 ( .A(N283), .B(N3063), .Y(N3286) );
  AND2X1 gate861 ( .A(N303), .B(N3064), .Y(N3287) );
  AND2X1 gate862 ( .A(N706), .B(N3065), .Y(N3288) );
  AND2X1 gate863 ( .A(N715), .B(N3066), .Y(N3289) );
  AND2X1 gate864 ( .A(N727), .B(N3067), .Y(N3290) );
  AND2X1 gate865 ( .A(N740), .B(N3068), .Y(N3291) );
  AND2X1 gate866 ( .A(N753), .B(N3069), .Y(N3292) );
  AND2X1 gate867 ( .A(N283), .B(N3070), .Y(N3293) );
  AND2X1 gate868 ( .A(N294), .B(N3071), .Y(N3294) );
  AND2X1 gate869 ( .A(N311), .B(N3072), .Y(N3295) );
  AND2X1 gate870 ( .A(N715), .B(N3073), .Y(N3296) );
  AND2X1 gate871 ( .A(N727), .B(N3074), .Y(N3297) );
  AND2X1 gate872 ( .A(N740), .B(N3075), .Y(N3298) );
  AND2X1 gate873 ( .A(N753), .B(N3076), .Y(N3299) );
  AND2X1 gate874 ( .A(N283), .B(N3077), .Y(N3300) );
  AND2X1 gate875 ( .A(N294), .B(N3078), .Y(N3301) );
  AND2X1 gate876 ( .A(N303), .B(N3079), .Y(N3302) );
  AND2X1 gate877 ( .A(N317), .B(N3080), .Y(N3303) );
  AND2X1 gate878 ( .A(N727), .B(N3081), .Y(N3304) );
  AND2X1 gate879 ( .A(N740), .B(N3082), .Y(N3305) );
  AND2X1 gate880 ( .A(N753), .B(N3083), .Y(N3306) );
  AND2X1 gate881 ( .A(N283), .B(N3084), .Y(N3307) );
  AND2X1 gate882 ( .A(N294), .B(N3085), .Y(N3308) );
  AND2X1 gate883 ( .A(N303), .B(N3086), .Y(N3309) );
  AND2X1 gate884 ( .A(N311), .B(N3087), .Y(N3310) );
  AND2X1 gate885 ( .A(N322), .B(N3088), .Y(N3311) );
  AND2X1 gate886 ( .A(N740), .B(N3089), .Y(N3312) );
  AND2X1 gate887 ( .A(N753), .B(N3090), .Y(N3313) );
  AND2X1 gate888 ( .A(N283), .B(N3091), .Y(N3314) );
  AND2X1 gate889 ( .A(N294), .B(N3092), .Y(N3315) );
  AND2X1 gate890 ( .A(N303), .B(N3093), .Y(N3316) );
  AND2X1 gate891 ( .A(N311), .B(N3094), .Y(N3317) );
  AND2X1 gate892 ( .A(N317), .B(N3095), .Y(N3318) );
  AND2X1 gate893 ( .A(N326), .B(N3096), .Y(N3319) );
  AND2X1 gate894 ( .A(N753), .B(N3097), .Y(N3320) );
  AND2X1 gate895 ( .A(N283), .B(N3098), .Y(N3321) );
  AND2X1 gate896 ( .A(N294), .B(N3099), .Y(N3322) );
  AND2X1 gate897 ( .A(N303), .B(N3100), .Y(N3323) );
  AND2X1 gate898 ( .A(N311), .B(N3101), .Y(N3324) );
  AND2X1 gate899 ( .A(N317), .B(N3102), .Y(N3325) );
  AND2X1 gate900 ( .A(N322), .B(N3103), .Y(N3326) );
  AND2X1 gate901 ( .A(N329), .B(N3104), .Y(N3327) );
  AND2X1 gate902 ( .A(N283), .B(N3105), .Y(N3328) );
  AND2X1 gate903 ( .A(N294), .B(N3106), .Y(N3329) );
  AND2X1 gate904 ( .A(N303), .B(N3107), .Y(N3330) );
  AND2X1 gate905 ( .A(N311), .B(N3108), .Y(N3331) );
  AND2X1 gate906 ( .A(N317), .B(N3109), .Y(N3332) );
  AND2X1 gate907 ( .A(N322), .B(N3110), .Y(N3333) );
  AND2X1 gate908 ( .A(N326), .B(N3111), .Y(N3334) );
  AND2X1 gate909_1 ( .A(N3190), .B(N3191), .Y(N3383_1) );
  AND2X1 gate909_2 ( .A(N3192), .B(N3193), .Y(N3383_2) );
  AND2X1 gate909_3 ( .A(N917), .B(N3383_1), .Y(N3383_3) );
  AND2X1 gate909 ( .A(N3383_2), .B(N3383_3), .Y(N3383) );
  BUFX2 gate910 ( .A(N2977), .Y(N3384) );
  AND2X1 gate911 ( .A(N3196), .B(N1736), .Y(N3387) );
  AND2X1 gate912 ( .A(N2977), .B(N2149), .Y(N3388) );
  AND2X1 gate913 ( .A(N2973), .B(N1737), .Y(N3389) );
  NOR3X1 gate914_1 ( .A(N3207), .B(N3208), .C(N3209), .Y(N3390_1) );
  NOR3X1 gate914_2 ( .A(N3210), .B(N3211), .C(N3212), .Y(N3390_2) );
  NOR3X1 gate914_3 ( .A(N3213), .B(N3214), .C(N3390_1), .Y(N3390_3) );
  NOR2X1 gate914 ( .A(N3390_2), .B(N3390_3), .Y(N3390) );
  NOR3X1 gate915_1 ( .A(N3215), .B(N3216), .C(N3217), .Y(N3391_1) );
  NOR3X1 gate915_2 ( .A(N3218), .B(N3219), .C(N3220), .Y(N3391_2) );
  NOR3X1 gate915_3 ( .A(N3221), .B(N3222), .C(N3391_1), .Y(N3391_3) );
  NOR2X1 gate915 ( .A(N3391_2), .B(N3391_3), .Y(N3391) );
  NOR3X1 gate916_1 ( .A(N3223), .B(N3224), .C(N3225), .Y(N3392_1) );
  NOR3X1 gate916_2 ( .A(N3226), .B(N3227), .C(N3228), .Y(N3392_2) );
  NOR3X1 gate916_3 ( .A(N3229), .B(N3230), .C(N3392_1), .Y(N3392_3) );
  NOR2X1 gate916 ( .A(N3392_2), .B(N3392_3), .Y(N3392) );
  NOR3X1 gate917_1 ( .A(N3231), .B(N3232), .C(N3233), .Y(N3393_1) );
  NOR3X1 gate917_2 ( .A(N3234), .B(N3235), .C(N3236), .Y(N3393_2) );
  NOR3X1 gate917_3 ( .A(N3237), .B(N3238), .C(N3393_1), .Y(N3393_3) );
  NOR2X1 gate917 ( .A(N3393_2), .B(N3393_3), .Y(N3393) );
  NOR3X1 gate918_1 ( .A(N3239), .B(N3240), .C(N3241), .Y(N3394_1) );
  NOR3X1 gate918_2 ( .A(N3242), .B(N3243), .C(N3244), .Y(N3394_2) );
  NOR3X1 gate918_3 ( .A(N3245), .B(N3246), .C(N3394_1), .Y(N3394_3) );
  NOR2X1 gate918 ( .A(N3394_2), .B(N3394_3), .Y(N3394) );
  NOR3X1 gate919_1 ( .A(N3247), .B(N3248), .C(N3249), .Y(N3395_1) );
  NOR3X1 gate919_2 ( .A(N3250), .B(N3251), .C(N3252), .Y(N3395_2) );
  NOR3X1 gate919_3 ( .A(N3253), .B(N3254), .C(N3395_1), .Y(N3395_3) );
  NOR2X1 gate919 ( .A(N3395_2), .B(N3395_3), .Y(N3395) );
  NOR3X1 gate920_1 ( .A(N3255), .B(N3256), .C(N3257), .Y(N3396_1) );
  NOR3X1 gate920_2 ( .A(N3258), .B(N3259), .C(N3260), .Y(N3396_2) );
  NOR3X1 gate920_3 ( .A(N3261), .B(N3262), .C(N3396_1), .Y(N3396_3) );
  NOR2X1 gate920 ( .A(N3396_2), .B(N3396_3), .Y(N3396) );
  NOR3X1 gate921_1 ( .A(N3263), .B(N3264), .C(N3265), .Y(N3397_1) );
  NOR3X1 gate921_2 ( .A(N3266), .B(N3267), .C(N3268), .Y(N3397_2) );
  NOR3X1 gate921_3 ( .A(N3269), .B(N3270), .C(N3397_1), .Y(N3397_3) );
  NOR2X1 gate921 ( .A(N3397_2), .B(N3397_3), .Y(N3397) );
  NOR3X1 gate922_1 ( .A(N3271), .B(N3272), .C(N3273), .Y(N3398_1) );
  NOR3X1 gate922_2 ( .A(N3274), .B(N3275), .C(N3276), .Y(N3398_2) );
  NOR3X1 gate922_3 ( .A(N3277), .B(N3278), .C(N3398_1), .Y(N3398_3) );
  NOR2X1 gate922 ( .A(N3398_2), .B(N3398_3), .Y(N3398) );
  NOR3X1 gate923_1 ( .A(N3279), .B(N3280), .C(N3281), .Y(N3399_1) );
  NOR3X1 gate923_2 ( .A(N3282), .B(N3283), .C(N3284), .Y(N3399_2) );
  NOR3X1 gate923_3 ( .A(N3285), .B(N3286), .C(N3399_1), .Y(N3399_3) );
  NOR2X1 gate923 ( .A(N3399_2), .B(N3399_3), .Y(N3399) );
  NOR3X1 gate924_1 ( .A(N3287), .B(N3288), .C(N3289), .Y(N3400_1) );
  NOR3X1 gate924_2 ( .A(N3290), .B(N3291), .C(N3292), .Y(N3400_2) );
  NOR3X1 gate924_3 ( .A(N3293), .B(N3294), .C(N3400_1), .Y(N3400_3) );
  NOR2X1 gate924 ( .A(N3400_2), .B(N3400_3), .Y(N3400) );
  NOR3X1 gate925_1 ( .A(N3295), .B(N3296), .C(N3297), .Y(N3401_1) );
  NOR3X1 gate925_2 ( .A(N3298), .B(N3299), .C(N3300), .Y(N3401_2) );
  NOR3X1 gate925_3 ( .A(N3301), .B(N3302), .C(N3401_1), .Y(N3401_3) );
  NOR2X1 gate925 ( .A(N3401_2), .B(N3401_3), .Y(N3401) );
  NOR3X1 gate926_1 ( .A(N3303), .B(N3304), .C(N3305), .Y(N3402_1) );
  NOR3X1 gate926_2 ( .A(N3306), .B(N3307), .C(N3308), .Y(N3402_2) );
  NOR3X1 gate926_3 ( .A(N3309), .B(N3310), .C(N3402_1), .Y(N3402_3) );
  NOR2X1 gate926 ( .A(N3402_2), .B(N3402_3), .Y(N3402) );
  NOR3X1 gate927_1 ( .A(N3311), .B(N3312), .C(N3313), .Y(N3403_1) );
  NOR3X1 gate927_2 ( .A(N3314), .B(N3315), .C(N3316), .Y(N3403_2) );
  NOR3X1 gate927_3 ( .A(N3317), .B(N3318), .C(N3403_1), .Y(N3403_3) );
  NOR2X1 gate927 ( .A(N3403_2), .B(N3403_3), .Y(N3403) );
  NOR3X1 gate928_1 ( .A(N3319), .B(N3320), .C(N3321), .Y(N3404_1) );
  NOR3X1 gate928_2 ( .A(N3322), .B(N3323), .C(N3324), .Y(N3404_2) );
  NOR3X1 gate928_3 ( .A(N3325), .B(N3326), .C(N3404_1), .Y(N3404_3) );
  NOR2X1 gate928 ( .A(N3404_2), .B(N3404_3), .Y(N3404) );
  NOR3X1 gate929_1 ( .A(N3327), .B(N3328), .C(N3329), .Y(N3405_1) );
  NOR3X1 gate929_2 ( .A(N3330), .B(N3331), .C(N3332), .Y(N3405_2) );
  NOR3X1 gate929_3 ( .A(N3333), .B(N3334), .C(N3405_1), .Y(N3405_3) );
  NOR2X1 gate929 ( .A(N3405_2), .B(N3405_3), .Y(N3405) );
  AND2X1 gate930 ( .A(N3206), .B(N2641), .Y(N3406) );
  AND2X1 gate931_1 ( .A(N169), .B(N2648), .Y(N3407_1) );
  AND2X1 gate931 ( .A(N3112), .B(N3407_1), .Y(N3407) );
  AND2X1 gate932_1 ( .A(N179), .B(N2648), .Y(N3410_1) );
  AND2X1 gate932 ( .A(N3115), .B(N3410_1), .Y(N3410) );
  AND2X1 gate933_1 ( .A(N190), .B(N2652), .Y(N3413_1) );
  AND2X1 gate933 ( .A(N3115), .B(N3413_1), .Y(N3413) );
  AND2X1 gate934_1 ( .A(N200), .B(N2652), .Y(N3414_1) );
  AND2X1 gate934 ( .A(N3112), .B(N3414_1), .Y(N3414) );
  OR2X1 gate935_1 ( .A(N3119), .B(N1875), .Y(N3415_1) );
  OR2X1 gate935 ( .A(N2073), .B(N3415_1), .Y(N3415) );
  NOR3X1 gate936 ( .A(N3119), .B(N1875), .C(N2073), .Y(N3419) );
  AND2X1 gate937_1 ( .A(N169), .B(N2662), .Y(N3423_1) );
  AND2X1 gate937 ( .A(N3128), .B(N3423_1), .Y(N3423) );
  AND2X1 gate938_1 ( .A(N179), .B(N2662), .Y(N3426_1) );
  AND2X1 gate938 ( .A(N3131), .B(N3426_1), .Y(N3426) );
  AND2X1 gate939_1 ( .A(N190), .B(N2666), .Y(N3429_1) );
  AND2X1 gate939 ( .A(N3131), .B(N3429_1), .Y(N3429) );
  AND2X1 gate940_1 ( .A(N200), .B(N2666), .Y(N3430_1) );
  AND2X1 gate940 ( .A(N3128), .B(N3430_1), .Y(N3430) );
  AND2X1 gate941_1 ( .A(N169), .B(N2673), .Y(N3431_1) );
  AND2X1 gate941 ( .A(N3135), .B(N3431_1), .Y(N3431) );
  AND2X1 gate942_1 ( .A(N179), .B(N2673), .Y(N3434_1) );
  AND2X1 gate942 ( .A(N3138), .B(N3434_1), .Y(N3434) );
  AND2X1 gate943_1 ( .A(N190), .B(N2677), .Y(N3437_1) );
  AND2X1 gate943 ( .A(N3138), .B(N3437_1), .Y(N3437) );
  AND2X1 gate944_1 ( .A(N200), .B(N2677), .Y(N3438_1) );
  AND2X1 gate944 ( .A(N3135), .B(N3438_1), .Y(N3438) );
  AND2X1 gate945_1 ( .A(N169), .B(N2684), .Y(N3439_1) );
  AND2X1 gate945 ( .A(N3142), .B(N3439_1), .Y(N3439) );
  AND2X1 gate946_1 ( .A(N179), .B(N2684), .Y(N3442_1) );
  AND2X1 gate946 ( .A(N3145), .B(N3442_1), .Y(N3442) );
  AND2X1 gate947_1 ( .A(N190), .B(N2688), .Y(N3445_1) );
  AND2X1 gate947 ( .A(N3145), .B(N3445_1), .Y(N3445) );
  AND2X1 gate948_1 ( .A(N200), .B(N2688), .Y(N3446_1) );
  AND2X1 gate948 ( .A(N3142), .B(N3446_1), .Y(N3446) );
  OR2X1 gate949_1 ( .A(N3149), .B(N1895), .Y(N3447_1) );
  OR2X1 gate949 ( .A(N2093), .B(N3447_1), .Y(N3447) );
  NOR3X1 gate950 ( .A(N3149), .B(N1895), .C(N2093), .Y(N3451) );
  AND2X1 gate951_1 ( .A(N169), .B(N2702), .Y(N3455_1) );
  AND2X1 gate951 ( .A(N3158), .B(N3455_1), .Y(N3455) );
  AND2X1 gate952_1 ( .A(N179), .B(N2702), .Y(N3458_1) );
  AND2X1 gate952 ( .A(N3161), .B(N3458_1), .Y(N3458) );
  AND2X1 gate953_1 ( .A(N190), .B(N2706), .Y(N3461_1) );
  AND2X1 gate953 ( .A(N3161), .B(N3461_1), .Y(N3461) );
  AND2X1 gate954_1 ( .A(N200), .B(N2706), .Y(N3462_1) );
  AND2X1 gate954 ( .A(N3158), .B(N3462_1), .Y(N3462) );
  AND2X1 gate955_1 ( .A(N169), .B(N2715), .Y(N3463_1) );
  AND2X1 gate955 ( .A(N3165), .B(N3463_1), .Y(N3463) );
  AND2X1 gate956_1 ( .A(N179), .B(N2715), .Y(N3466_1) );
  AND2X1 gate956 ( .A(N3168), .B(N3466_1), .Y(N3466) );
  AND2X1 gate957_1 ( .A(N190), .B(N2719), .Y(N3469_1) );
  AND2X1 gate957 ( .A(N3168), .B(N3469_1), .Y(N3469) );
  AND2X1 gate958_1 ( .A(N200), .B(N2719), .Y(N3470_1) );
  AND2X1 gate958 ( .A(N3165), .B(N3470_1), .Y(N3470) );
  OR2X1 gate959 ( .A(N3194), .B(N3383), .Y(N3471) );
  BUFX2 gate960 ( .A(N2967), .Y(N3472) );
  BUFX2 gate961 ( .A(N2970), .Y(N3475) );
  BUFX2 gate962 ( .A(N2967), .Y(N3478) );
  BUFX2 gate963 ( .A(N2970), .Y(N3481) );
  BUFX2 gate964 ( .A(N2973), .Y(N3484) );
  BUFX2 gate965 ( .A(N2973), .Y(N3487) );
  BUFX2 gate966 ( .A(N3172), .Y(N3490) );
  BUFX2 gate967 ( .A(N3172), .Y(N3493) );
  BUFX2 gate968 ( .A(N3175), .Y(N3496) );
  BUFX2 gate969 ( .A(N3175), .Y(N3499) );
  BUFX2 gate970 ( .A(N3178), .Y(N3502) );
  BUFX2 gate971 ( .A(N3178), .Y(N3505) );
  BUFX2 gate972 ( .A(N3181), .Y(N3508) );
  BUFX2 gate973 ( .A(N3181), .Y(N3511) );
  BUFX2 gate974 ( .A(N3184), .Y(N3514) );
  BUFX2 gate975 ( .A(N3184), .Y(N3517) );
  BUFX2 gate976 ( .A(N3187), .Y(N3520) );
  BUFX2 gate977 ( .A(N3187), .Y(N3523) );
  NOR2X1 gate978 ( .A(N3387), .B(N2350), .Y(N3534) );
  OR2X1 gate979_1 ( .A(N3388), .B(N2151), .Y(N3535_1) );
  OR2X1 gate979 ( .A(N2351), .B(N3535_1), .Y(N3535) );
  NOR2X1 gate980 ( .A(N3389), .B(N1966), .Y(N3536) );
  AND2X1 gate981 ( .A(N3390), .B(N2209), .Y(N3537) );
  AND2X1 gate982 ( .A(N3398), .B(N2210), .Y(N3538) );
  AND2X1 gate983 ( .A(N3391), .B(N1842), .Y(N3539) );
  AND2X1 gate984 ( .A(N3399), .B(N1369), .Y(N3540) );
  AND2X1 gate985 ( .A(N3392), .B(N1843), .Y(N3541) );
  AND2X1 gate986 ( .A(N3400), .B(N1369), .Y(N3542) );
  AND2X1 gate987 ( .A(N3393), .B(N1844), .Y(N3543) );
  AND2X1 gate988 ( .A(N3401), .B(N1369), .Y(N3544) );
  AND2X1 gate989 ( .A(N3394), .B(N1845), .Y(N3545) );
  AND2X1 gate990 ( .A(N3402), .B(N1369), .Y(N3546) );
  AND2X1 gate991 ( .A(N3395), .B(N1846), .Y(N3547) );
  AND2X1 gate992 ( .A(N3403), .B(N1369), .Y(N3548) );
  AND2X1 gate993 ( .A(N3396), .B(N1847), .Y(N3549) );
  AND2X1 gate994 ( .A(N3404), .B(N1369), .Y(N3550) );
  AND2X1 gate995 ( .A(N3397), .B(N1848), .Y(N3551) );
  AND2X1 gate996 ( .A(N3405), .B(N1369), .Y(N3552) );
  OR2X1 gate997_1 ( .A(N3413), .B(N3414), .Y(N3557_1) );
  OR2X1 gate997 ( .A(N3118), .B(N3557_1), .Y(N3557) );
  OR2X1 gate998_1 ( .A(N3429), .B(N3430), .Y(N3568_1) );
  OR2X1 gate998 ( .A(N3134), .B(N3568_1), .Y(N3568) );
  OR2X1 gate999_1 ( .A(N3437), .B(N3438), .Y(N3573_1) );
  OR2X1 gate999 ( .A(N3141), .B(N3573_1), .Y(N3573) );
  OR2X1 gate1000_1 ( .A(N3445), .B(N3446), .Y(N3578_1) );
  OR2X1 gate1000 ( .A(N3148), .B(N3578_1), .Y(N3578) );
  OR2X1 gate1001_1 ( .A(N3461), .B(N3462), .Y(N3589_1) );
  OR2X1 gate1001 ( .A(N3164), .B(N3589_1), .Y(N3589) );
  OR2X1 gate1002_1 ( .A(N3469), .B(N3470), .Y(N3594_1) );
  OR2X1 gate1002 ( .A(N3171), .B(N3594_1), .Y(N3594) );
  AND2X1 gate1003 ( .A(N3471), .B(N2728), .Y(N3605) );
  INVX1 gate1004 ( .A(N3478), .Y(N3626) );
  INVX1 gate1005 ( .A(N3481), .Y(N3627) );
  INVX1 gate1006 ( .A(N3487), .Y(N3628) );
  INVX1 gate1007 ( .A(N3484), .Y(N3629) );
  INVX1 gate1008 ( .A(N3472), .Y(N3630) );
  INVX1 gate1009 ( .A(N3475), .Y(N3631) );
  AND2X1 gate1010 ( .A(N3536), .B(N2152), .Y(N3632) );
  AND2X1 gate1011 ( .A(N3534), .B(N2155), .Y(N3633) );
  OR2X1 gate1012_1 ( .A(N3537), .B(N3538), .Y(N3634_1) );
  OR2X1 gate1012 ( .A(N2398), .B(N3634_1), .Y(N3634) );
  OR2X1 gate1013 ( .A(N3539), .B(N3540), .Y(N3635) );
  OR2X1 gate1014 ( .A(N3541), .B(N3542), .Y(N3636) );
  OR2X1 gate1015 ( .A(N3543), .B(N3544), .Y(N3637) );
  OR2X1 gate1016 ( .A(N3545), .B(N3546), .Y(N3638) );
  OR2X1 gate1017 ( .A(N3547), .B(N3548), .Y(N3639) );
  OR2X1 gate1018 ( .A(N3549), .B(N3550), .Y(N3640) );
  OR2X1 gate1019 ( .A(N3551), .B(N3552), .Y(N3641) );
  AND2X1 gate1020 ( .A(N3535), .B(N2643), .Y(N3642) );
  OR2X1 gate1021 ( .A(N3407), .B(N3410), .Y(N3643) );
  NOR2X1 gate1022 ( .A(N3407), .B(N3410), .Y(N3644) );
  AND2X1 gate1023_1 ( .A(N169), .B(N3415), .Y(N3645_1) );
  AND2X1 gate1023 ( .A(N3122), .B(N3645_1), .Y(N3645) );
  AND2X1 gate1024_1 ( .A(N179), .B(N3415), .Y(N3648_1) );
  AND2X1 gate1024 ( .A(N3125), .B(N3648_1), .Y(N3648) );
  AND2X1 gate1025_1 ( .A(N190), .B(N3419), .Y(N3651_1) );
  AND2X1 gate1025 ( .A(N3125), .B(N3651_1), .Y(N3651) );
  AND2X1 gate1026_1 ( .A(N200), .B(N3419), .Y(N3652_1) );
  AND2X1 gate1026 ( .A(N3122), .B(N3652_1), .Y(N3652) );
  INVX1 gate1027 ( .A(N3419), .Y(N3653) );
  OR2X1 gate1028 ( .A(N3423), .B(N3426), .Y(N3654) );
  NOR2X1 gate1029 ( .A(N3423), .B(N3426), .Y(N3657) );
  OR2X1 gate1030 ( .A(N3431), .B(N3434), .Y(N3658) );
  NOR2X1 gate1031 ( .A(N3431), .B(N3434), .Y(N3661) );
  OR2X1 gate1032 ( .A(N3439), .B(N3442), .Y(N3662) );
  NOR2X1 gate1033 ( .A(N3439), .B(N3442), .Y(N3663) );
  AND2X1 gate1034_1 ( .A(N169), .B(N3447), .Y(N3664_1) );
  AND2X1 gate1034 ( .A(N3152), .B(N3664_1), .Y(N3664) );
  AND2X1 gate1035_1 ( .A(N179), .B(N3447), .Y(N3667_1) );
  AND2X1 gate1035 ( .A(N3155), .B(N3667_1), .Y(N3667) );
  AND2X1 gate1036_1 ( .A(N190), .B(N3451), .Y(N3670_1) );
  AND2X1 gate1036 ( .A(N3155), .B(N3670_1), .Y(N3670) );
  AND2X1 gate1037_1 ( .A(N200), .B(N3451), .Y(N3671_1) );
  AND2X1 gate1037 ( .A(N3152), .B(N3671_1), .Y(N3671) );
  INVX1 gate1038 ( .A(N3451), .Y(N3672) );
  OR2X1 gate1039 ( .A(N3455), .B(N3458), .Y(N3673) );
  NOR2X1 gate1040 ( .A(N3455), .B(N3458), .Y(N3676) );
  OR2X1 gate1041 ( .A(N3463), .B(N3466), .Y(N3677) );
  NOR2X1 gate1042 ( .A(N3463), .B(N3466), .Y(N3680) );
  INVX1 gate1043 ( .A(N3493), .Y(N3681) );
  AND2X1 gate1044 ( .A(N1909), .B(N3415), .Y(N3682) );
  INVX1 gate1045 ( .A(N3496), .Y(N3685) );
  INVX1 gate1046 ( .A(N3499), .Y(N3686) );
  INVX1 gate1047 ( .A(N3502), .Y(N3687) );
  INVX1 gate1048 ( .A(N3505), .Y(N3688) );
  INVX1 gate1049 ( .A(N3511), .Y(N3689) );
  AND2X1 gate1050 ( .A(N1922), .B(N3447), .Y(N3690) );
  INVX1 gate1051 ( .A(N3517), .Y(N3693) );
  INVX1 gate1052 ( .A(N3520), .Y(N3694) );
  INVX1 gate1053 ( .A(N3523), .Y(N3695) );
  INVX1 gate1054 ( .A(N3514), .Y(N3696) );
  BUFX2 gate1055 ( .A(N3384), .Y(N3697) );
  BUFX2 gate1056 ( .A(N3384), .Y(N3700) );
  INVX1 gate1057 ( .A(N3490), .Y(N3703) );
  INVX1 gate1058 ( .A(N3508), .Y(N3704) );
  NAND2X1 gate1059 ( .A(N3475), .B(N3630), .Y(N3705) );
  NAND2X1 gate1060 ( .A(N3472), .B(N3631), .Y(N3706) );
  NAND2X1 gate1061 ( .A(N3481), .B(N3626), .Y(N3707) );
  NAND2X1 gate1062 ( .A(N3478), .B(N3627), .Y(N3708) );
  OR2X1 gate1063_1 ( .A(N3632), .B(N2352), .Y(N3711_1) );
  OR2X1 gate1063 ( .A(N2353), .B(N3711_1), .Y(N3711) );
  OR2X1 gate1064_1 ( .A(N3633), .B(N2354), .Y(N3712_1) );
  OR2X1 gate1064 ( .A(N2355), .B(N3712_1), .Y(N3712) );
  AND2X1 gate1065 ( .A(N3634), .B(N2632), .Y(N3713) );
  AND2X1 gate1066 ( .A(N3635), .B(N2634), .Y(N3714) );
  AND2X1 gate1067 ( .A(N3636), .B(N2636), .Y(N3715) );
  AND2X1 gate1068 ( .A(N3637), .B(N2638), .Y(N3716) );
  AND2X1 gate1069 ( .A(N3638), .B(N2640), .Y(N3717) );
  AND2X1 gate1070 ( .A(N3639), .B(N2642), .Y(N3718) );
  AND2X1 gate1071 ( .A(N3640), .B(N2644), .Y(N3719) );
  AND2X1 gate1072 ( .A(N3641), .B(N2646), .Y(N3720) );
  AND2X1 gate1073 ( .A(N3644), .B(N3557), .Y(N3721) );
  OR2X1 gate1074_1 ( .A(N3651), .B(N3652), .Y(N3731_1) );
  OR2X1 gate1074 ( .A(N3653), .B(N3731_1), .Y(N3731) );
  AND2X1 gate1075 ( .A(N3657), .B(N3568), .Y(N3734) );
  AND2X1 gate1076 ( .A(N3661), .B(N3573), .Y(N3740) );
  AND2X1 gate1077 ( .A(N3663), .B(N3578), .Y(N3743) );
  OR2X1 gate1078_1 ( .A(N3670), .B(N3671), .Y(N3753_1) );
  OR2X1 gate1078 ( .A(N3672), .B(N3753_1), .Y(N3753) );
  AND2X1 gate1079 ( .A(N3676), .B(N3589), .Y(N3756) );
  AND2X1 gate1080 ( .A(N3680), .B(N3594), .Y(N3762) );
  INVX1 gate1081 ( .A(N3643), .Y(N3765) );
  INVX1 gate1082 ( .A(N3662), .Y(N3766) );
  NAND2X1 gate1083 ( .A(N3705), .B(N3706), .Y(N3773) );
  NAND2X1 gate1084 ( .A(N3707), .B(N3708), .Y(N3774) );
  NAND2X1 gate1085 ( .A(N3700), .B(N3628), .Y(N3775) );
  INVX1 gate1086 ( .A(N3700), .Y(N3776) );
  NAND2X1 gate1087 ( .A(N3697), .B(N3629), .Y(N3777) );
  INVX1 gate1088 ( .A(N3697), .Y(N3778) );
  AND2X1 gate1089 ( .A(N3712), .B(N2645), .Y(N3779) );
  AND2X1 gate1090 ( .A(N3711), .B(N2647), .Y(N3780) );
  OR2X1 gate1091 ( .A(N3645), .B(N3648), .Y(N3786) );
  NOR2X1 gate1092 ( .A(N3645), .B(N3648), .Y(N3789) );
  OR2X1 gate1093 ( .A(N3664), .B(N3667), .Y(N3800) );
  NOR2X1 gate1094 ( .A(N3664), .B(N3667), .Y(N3803) );
  AND2X1 gate1095 ( .A(N3654), .B(N1917), .Y(N3809) );
  AND2X1 gate1096 ( .A(N3658), .B(N1917), .Y(N3812) );
  AND2X1 gate1097 ( .A(N3673), .B(N1926), .Y(N3815) );
  AND2X1 gate1098 ( .A(N3677), .B(N1926), .Y(N3818) );
  BUFX2 gate1099 ( .A(N3682), .Y(N3821) );
  BUFX2 gate1100 ( .A(N3682), .Y(N3824) );
  BUFX2 gate1101 ( .A(N3690), .Y(N3827) );
  BUFX2 gate1102 ( .A(N3690), .Y(N3830) );
  NAND2X1 gate1103 ( .A(N3773), .B(N3774), .Y(N3833) );
  NAND2X1 gate1104 ( .A(N3487), .B(N3776), .Y(N3834) );
  NAND2X1 gate1105 ( .A(N3484), .B(N3778), .Y(N3835) );
  AND2X1 gate1106 ( .A(N3789), .B(N3731), .Y(N3838) );
  AND2X1 gate1107 ( .A(N3803), .B(N3753), .Y(N3845) );
  BUFX2 gate1108 ( .A(N3721), .Y(N3850) );
  BUFX2 gate1109 ( .A(N3734), .Y(N3855) );
  BUFX2 gate1110 ( .A(N3740), .Y(N3858) );
  BUFX2 gate1111 ( .A(N3743), .Y(N3861) );
  BUFX2 gate1112 ( .A(N3756), .Y(N3865) );
  BUFX2 gate1113 ( .A(N3762), .Y(N3868) );
  NAND2X1 gate1114 ( .A(N3775), .B(N3834), .Y(N3884) );
  NAND2X1 gate1115 ( .A(N3777), .B(N3835), .Y(N3885) );
  NAND2X1 gate1116 ( .A(N3721), .B(N3786), .Y(N3894) );
  NAND2X1 gate1117 ( .A(N3743), .B(N3800), .Y(N3895) );
  INVX1 gate1118 ( .A(N3821), .Y(N3898) );
  INVX1 gate1119 ( .A(N3824), .Y(N3899) );
  INVX1 gate1120 ( .A(N3830), .Y(N3906) );
  INVX1 gate1121 ( .A(N3827), .Y(N3911) );
  AND2X1 gate1122 ( .A(N3786), .B(N1912), .Y(N3912) );
  BUFX2 gate1123 ( .A(N3812), .Y(N3913) );
  AND2X1 gate1124 ( .A(N3800), .B(N1917), .Y(N3916) );
  BUFX2 gate1125 ( .A(N3818), .Y(N3917) );
  INVX1 gate1126 ( .A(N3809), .Y(N3920) );
  BUFX2 gate1127 ( .A(N3818), .Y(N3921) );
  INVX1 gate1128 ( .A(N3884), .Y(N3924) );
  INVX1 gate1129 ( .A(N3885), .Y(N3925) );
  AND2X1 gate1130_1 ( .A(N3721), .B(N3838), .Y(N3926_1) );
  AND2X1 gate1130_2 ( .A(N3734), .B(N3740), .Y(N3926_2) );
  AND2X1 gate1130 ( .A(N3926_1), .B(N3926_2), .Y(N3926) );
  NAND3X1 gate1131 ( .A(N3721), .B(N3838), .C(N3654), .Y(N3930) );
  NAND2X1 gate1132_1 ( .A(N3658), .B(N3838), .Y(N3931_1) );
  NAND2X1 gate1132_2 ( .A(N3734), .B(N3721), .Y(N3931_2) );
  NAND2X1 gate1132 ( .A(N3931_1), .B(N3931_2), .Y(N3931) );
  AND2X1 gate1133_1 ( .A(N3743), .B(N3845), .Y(N3932_1) );
  AND2X1 gate1133_2 ( .A(N3756), .B(N3762), .Y(N3932_2) );
  AND2X1 gate1133 ( .A(N3932_1), .B(N3932_2), .Y(N3932) );
  NAND3X1 gate1134 ( .A(N3743), .B(N3845), .C(N3673), .Y(N3935) );
  NAND2X1 gate1135_1 ( .A(N3677), .B(N3845), .Y(N3936_1) );
  NAND2X1 gate1135_2 ( .A(N3756), .B(N3743), .Y(N3936_2) );
  NAND2X1 gate1135 ( .A(N3936_1), .B(N3936_2), .Y(N3936) );
  BUFX2 gate1136 ( .A(N3838), .Y(N3937) );
  BUFX2 gate1137 ( .A(N3845), .Y(N3940) );
  INVX1 gate1138 ( .A(N3912), .Y(N3947) );
  INVX1 gate1139 ( .A(N3916), .Y(N3948) );
  BUFX2 gate1140 ( .A(N3850), .Y(N3950) );
  BUFX2 gate1141 ( .A(N3850), .Y(N3953) );
  BUFX2 gate1142 ( .A(N3855), .Y(N3956) );
  BUFX2 gate1143 ( .A(N3855), .Y(N3959) );
  BUFX2 gate1144 ( .A(N3858), .Y(N3962) );
  BUFX2 gate1145 ( .A(N3858), .Y(N3965) );
  BUFX2 gate1146 ( .A(N3861), .Y(N3968) );
  BUFX2 gate1147 ( .A(N3861), .Y(N3971) );
  BUFX2 gate1148 ( .A(N3865), .Y(N3974) );
  BUFX2 gate1149 ( .A(N3865), .Y(N3977) );
  BUFX2 gate1150 ( .A(N3868), .Y(N3980) );
  BUFX2 gate1151 ( .A(N3868), .Y(N3983) );
  NAND2X1 gate1152 ( .A(N3924), .B(N3925), .Y(N3987) );
  NAND2X1 gate1153_1 ( .A(N3765), .B(N3894), .Y(N3992_1) );
  NAND2X1 gate1153_2 ( .A(N3930), .B(N3931), .Y(N3992_2) );
  NAND2X1 gate1153 ( .A(N3992_1), .B(N3992_2), .Y(N3992) );
  NAND2X1 gate1154_1 ( .A(N3766), .B(N3895), .Y(N3996_1) );
  NAND2X1 gate1154_2 ( .A(N3935), .B(N3936), .Y(N3996_2) );
  NAND2X1 gate1154 ( .A(N3996_1), .B(N3996_2), .Y(N3996) );
  INVX1 gate1155 ( .A(N3921), .Y(N4013) );
  AND2X1 gate1156 ( .A(N3932), .B(N3926), .Y(N4028) );
  NAND2X1 gate1157 ( .A(N3953), .B(N3681), .Y(N4029) );
  NAND2X1 gate1158 ( .A(N3959), .B(N3686), .Y(N4030) );
  NAND2X1 gate1159 ( .A(N3965), .B(N3688), .Y(N4031) );
  NAND2X1 gate1160 ( .A(N3971), .B(N3689), .Y(N4032) );
  NAND2X1 gate1161 ( .A(N3977), .B(N3693), .Y(N4033) );
  NAND2X1 gate1162 ( .A(N3983), .B(N3695), .Y(N4034) );
  BUFX2 gate1163 ( .A(N3926), .Y(N4035) );
  INVX1 gate1164 ( .A(N3953), .Y(N4042) );
  INVX1 gate1165 ( .A(N3956), .Y(N4043) );
  NAND2X1 gate1166 ( .A(N3956), .B(N3685), .Y(N4044) );
  INVX1 gate1167 ( .A(N3959), .Y(N4045) );
  INVX1 gate1168 ( .A(N3962), .Y(N4046) );
  NAND2X1 gate1169 ( .A(N3962), .B(N3687), .Y(N4047) );
  INVX1 gate1170 ( .A(N3965), .Y(N4048) );
  INVX1 gate1171 ( .A(N3971), .Y(N4049) );
  INVX1 gate1172 ( .A(N3977), .Y(N4050) );
  INVX1 gate1173 ( .A(N3980), .Y(N4051) );
  NAND2X1 gate1174 ( .A(N3980), .B(N3694), .Y(N4052) );
  INVX1 gate1175 ( .A(N3983), .Y(N4053) );
  INVX1 gate1176 ( .A(N3974), .Y(N4054) );
  NAND2X1 gate1177 ( .A(N3974), .B(N3696), .Y(N4055) );
  AND2X1 gate1178 ( .A(N3932), .B(N2304), .Y(N4056) );
  INVX1 gate1179 ( .A(N3950), .Y(N4057) );
  NAND2X1 gate1180 ( .A(N3950), .B(N3703), .Y(N4058) );
  BUFX2 gate1181 ( .A(N3937), .Y(N4059) );
  BUFX2 gate1182 ( .A(N3937), .Y(N4062) );
  INVX1 gate1183 ( .A(N3968), .Y(N4065) );
  NAND2X1 gate1184 ( .A(N3968), .B(N3704), .Y(N4066) );
  BUFX2 gate1185 ( .A(N3940), .Y(N4067) );
  BUFX2 gate1186 ( .A(N3940), .Y(N4070) );
  NAND2X1 gate1187 ( .A(N3926), .B(N3996), .Y(N4073) );
  INVX1 gate1188 ( .A(N3992), .Y(N4074) );
  NAND2X1 gate1189 ( .A(N3493), .B(N4042), .Y(N4075) );
  NAND2X1 gate1190 ( .A(N3499), .B(N4045), .Y(N4076) );
  NAND2X1 gate1191 ( .A(N3505), .B(N4048), .Y(N4077) );
  NAND2X1 gate1192 ( .A(N3511), .B(N4049), .Y(N4078) );
  NAND2X1 gate1193 ( .A(N3517), .B(N4050), .Y(N4079) );
  NAND2X1 gate1194 ( .A(N3523), .B(N4053), .Y(N4080) );
  NAND2X1 gate1195 ( .A(N3496), .B(N4043), .Y(N4085) );
  NAND2X1 gate1196 ( .A(N3502), .B(N4046), .Y(N4086) );
  NAND2X1 gate1197 ( .A(N3520), .B(N4051), .Y(N4088) );
  NAND2X1 gate1198 ( .A(N3514), .B(N4054), .Y(N4090) );
  AND2X1 gate1199 ( .A(N3996), .B(N1926), .Y(N4091) );
  OR2X1 gate1200 ( .A(N3605), .B(N4056), .Y(N4094) );
  NAND2X1 gate1201 ( .A(N3490), .B(N4057), .Y(N4098) );
  NAND2X1 gate1202 ( .A(N3508), .B(N4065), .Y(N4101) );
  AND2X1 gate1203 ( .A(N4073), .B(N4074), .Y(N4104) );
  NAND2X1 gate1204 ( .A(N4075), .B(N4029), .Y(N4105) );
  NAND2X1 gate1205 ( .A(N4062), .B(N3899), .Y(N4106) );
  NAND2X1 gate1206 ( .A(N4076), .B(N4030), .Y(N4107) );
  NAND2X1 gate1207 ( .A(N4077), .B(N4031), .Y(N4108) );
  NAND2X1 gate1208 ( .A(N4078), .B(N4032), .Y(N4109) );
  NAND2X1 gate1209 ( .A(N4070), .B(N3906), .Y(N4110) );
  NAND2X1 gate1210 ( .A(N4079), .B(N4033), .Y(N4111) );
  NAND2X1 gate1211 ( .A(N4080), .B(N4034), .Y(N4112) );
  INVX1 gate1212 ( .A(N4059), .Y(N4113) );
  NAND2X1 gate1213 ( .A(N4059), .B(N3898), .Y(N4114) );
  INVX1 gate1214 ( .A(N4062), .Y(N4115) );
  NAND2X1 gate1215 ( .A(N4085), .B(N4044), .Y(N4116) );
  NAND2X1 gate1216 ( .A(N4086), .B(N4047), .Y(N4119) );
  INVX1 gate1217 ( .A(N4070), .Y(N4122) );
  NAND2X1 gate1218 ( .A(N4088), .B(N4052), .Y(N4123) );
  INVX1 gate1219 ( .A(N4067), .Y(N4126) );
  NAND2X1 gate1220 ( .A(N4067), .B(N3911), .Y(N4127) );
  NAND2X1 gate1221 ( .A(N4090), .B(N4055), .Y(N4128) );
  NAND2X1 gate1222 ( .A(N4098), .B(N4058), .Y(N4139) );
  NAND2X1 gate1223 ( .A(N4101), .B(N4066), .Y(N4142) );
  INVX1 gate1224 ( .A(N4104), .Y(N4145) );
  INVX1 gate1225 ( .A(N4105), .Y(N4146) );
  NAND2X1 gate1226 ( .A(N3824), .B(N4115), .Y(N4147) );
  INVX1 gate1227 ( .A(N4107), .Y(N4148) );
  INVX1 gate1228 ( .A(N4108), .Y(N4149) );
  INVX1 gate1229 ( .A(N4109), .Y(N4150) );
  NAND2X1 gate1230 ( .A(N3830), .B(N4122), .Y(N4151) );
  INVX1 gate1231 ( .A(N4111), .Y(N4152) );
  INVX1 gate1232 ( .A(N4112), .Y(N4153) );
  NAND2X1 gate1233 ( .A(N3821), .B(N4113), .Y(N4154) );
  NAND2X1 gate1234 ( .A(N3827), .B(N4126), .Y(N4161) );
  BUFX2 gate1235 ( .A(N4091), .Y(N4167) );
  BUFX2 gate1236 ( .A(N4094), .Y(N4174) );
  BUFX2 gate1237 ( .A(N4091), .Y(N4182) );
  AND2X1 gate1238 ( .A(N330), .B(N4094), .Y(N4186) );
  AND2X1 gate1239 ( .A(N4146), .B(N2230), .Y(N4189) );
  NAND2X1 gate1240 ( .A(N4147), .B(N4106), .Y(N4190) );
  AND2X1 gate1241 ( .A(N4148), .B(N2232), .Y(N4191) );
  AND2X1 gate1242 ( .A(N4149), .B(N2233), .Y(N4192) );
  AND2X1 gate1243 ( .A(N4150), .B(N2234), .Y(N4193) );
  NAND2X1 gate1244 ( .A(N4151), .B(N4110), .Y(N4194) );
  AND2X1 gate1245 ( .A(N4152), .B(N2236), .Y(N4195) );
  AND2X1 gate1246 ( .A(N4153), .B(N2237), .Y(N4196) );
  NAND2X1 gate1247 ( .A(N4154), .B(N4114), .Y(N4197) );
  BUFX2 gate1248 ( .A(N4116), .Y(N4200) );
  BUFX2 gate1249 ( .A(N4116), .Y(N4203) );
  BUFX2 gate1250 ( .A(N4119), .Y(N4209) );
  BUFX2 gate1251 ( .A(N4119), .Y(N4213) );
  NAND2X1 gate1252 ( .A(N4161), .B(N4127), .Y(N4218) );
  BUFX2 gate1253 ( .A(N4123), .Y(N4223) );
  AND2X1 gate1254 ( .A(N4128), .B(N3917), .Y(N4238) );
  INVX1 gate1255 ( .A(N4139), .Y(N4239) );
  INVX1 gate1256 ( .A(N4142), .Y(N4241) );
  AND2X1 gate1257 ( .A(N330), .B(N4123), .Y(N4242) );
  BUFX2 gate1258 ( .A(N4128), .Y(N4247) );
  NOR3X1 gate1259 ( .A(N3713), .B(N4189), .C(N2898), .Y(N4251) );
  INVX1 gate1260 ( .A(N4190), .Y(N4252) );
  NOR3X1 gate1261 ( .A(N3715), .B(N4191), .C(N2900), .Y(N4253) );
  NOR3X1 gate1262 ( .A(N3716), .B(N4192), .C(N2901), .Y(N4254) );
  NOR3X1 gate1263 ( .A(N3717), .B(N4193), .C(N3406), .Y(N4255) );
  INVX1 gate1264 ( .A(N4194), .Y(N4256) );
  NOR3X1 gate1265 ( .A(N3719), .B(N4195), .C(N3779), .Y(N4257) );
  NOR3X1 gate1266 ( .A(N3720), .B(N4196), .C(N3780), .Y(N4258) );
  AND2X1 gate1267 ( .A(N4167), .B(N4035), .Y(N4283) );
  AND2X1 gate1268 ( .A(N4174), .B(N4035), .Y(N4284) );
  OR2X1 gate1269 ( .A(N3815), .B(N4238), .Y(N4287) );
  INVX1 gate1270 ( .A(N4186), .Y(N4291) );
  INVX1 gate1271 ( .A(N4167), .Y(N4295) );
  BUFX2 gate1272 ( .A(N4167), .Y(N4296) );
  INVX1 gate1273 ( .A(N4182), .Y(N4299) );
  AND2X1 gate1274 ( .A(N4252), .B(N2231), .Y(N4303) );
  AND2X1 gate1275 ( .A(N4256), .B(N2235), .Y(N4304) );
  BUFX2 gate1276 ( .A(N4197), .Y(N4305) );
  OR2X1 gate1277 ( .A(N3992), .B(N4283), .Y(N4310) );
  AND2X1 gate1278_1 ( .A(N4174), .B(N4213), .Y(N4316_1) );
  AND2X1 gate1278 ( .A(N4203), .B(N4316_1), .Y(N4316) );
  AND2X1 gate1279 ( .A(N4174), .B(N4209), .Y(N4317) );
  AND2X1 gate1280_1 ( .A(N4223), .B(N4128), .Y(N4318_1) );
  AND2X1 gate1280 ( .A(N4218), .B(N4318_1), .Y(N4318) );
  AND2X1 gate1281 ( .A(N4223), .B(N4128), .Y(N4319) );
  AND2X1 gate1282 ( .A(N4167), .B(N4209), .Y(N4322) );
  NAND2X1 gate1283 ( .A(N4203), .B(N3913), .Y(N4325) );
  NAND3X1 gate1284 ( .A(N4203), .B(N4213), .C(N4167), .Y(N4326) );
  NAND2X1 gate1285 ( .A(N4218), .B(N3815), .Y(N4327) );
  NAND3X1 gate1286 ( .A(N4218), .B(N4128), .C(N3917), .Y(N4328) );
  NAND2X1 gate1287 ( .A(N4247), .B(N4013), .Y(N4329) );
  INVX1 gate1288 ( .A(N4247), .Y(N4330) );
  AND2X1 gate1289_1 ( .A(N330), .B(N4094), .Y(N4331_1) );
  AND2X1 gate1289 ( .A(N4295), .B(N4331_1), .Y(N4331) );
  AND2X1 gate1290 ( .A(N4251), .B(N2730), .Y(N4335) );
  AND2X1 gate1291 ( .A(N4253), .B(N2734), .Y(N4338) );
  AND2X1 gate1292 ( .A(N4254), .B(N2736), .Y(N4341) );
  AND2X1 gate1293 ( .A(N4255), .B(N2738), .Y(N4344) );
  AND2X1 gate1294 ( .A(N4257), .B(N2742), .Y(N4347) );
  AND2X1 gate1295 ( .A(N4258), .B(N2744), .Y(N4350) );
  BUFX2 gate1296 ( .A(N4197), .Y(N4353) );
  BUFX2 gate1297 ( .A(N4203), .Y(N4356) );
  BUFX2 gate1298 ( .A(N4209), .Y(N4359) );
  BUFX2 gate1299 ( .A(N4218), .Y(N4362) );
  BUFX2 gate1300 ( .A(N4242), .Y(N4365) );
  BUFX2 gate1301 ( .A(N4242), .Y(N4368) );
  AND2X1 gate1302 ( .A(N4223), .B(N4223), .Y(N4371) );
  NOR3X1 gate1303 ( .A(N3714), .B(N4303), .C(N2899), .Y(N4376) );
  NOR3X1 gate1304 ( .A(N3718), .B(N4304), .C(N3642), .Y(N4377) );
  AND2X1 gate1305 ( .A(N330), .B(N4317), .Y(N4387) );
  AND2X1 gate1306 ( .A(N330), .B(N4318), .Y(N4390) );
  NAND2X1 gate1307 ( .A(N3921), .B(N4330), .Y(N4393) );
  BUFX2 gate1308 ( .A(N4287), .Y(N4398) );
  BUFX2 gate1309 ( .A(N4284), .Y(N4413) );
  NAND3X1 gate1310 ( .A(N3920), .B(N4325), .C(N4326), .Y(N4416) );
  OR2X1 gate1311 ( .A(N3812), .B(N4322), .Y(N4421) );
  NAND3X1 gate1312 ( .A(N3948), .B(N4327), .C(N4328), .Y(N4427) );
  BUFX2 gate1313 ( .A(N4287), .Y(N4430) );
  AND2X1 gate1314 ( .A(N330), .B(N4316), .Y(N4435) );
  OR2X1 gate1315 ( .A(N4331), .B(N4296), .Y(N4442) );
  AND2X1 gate1316_1 ( .A(N4174), .B(N4305), .Y(N4443_1) );
  AND2X1 gate1316_2 ( .A(N4203), .B(N4213), .Y(N4443_2) );
  AND2X1 gate1316 ( .A(N4443_1), .B(N4443_2), .Y(N4443) );
  NAND2X1 gate1317 ( .A(N4305), .B(N3809), .Y(N4446) );
  NAND3X1 gate1318 ( .A(N4305), .B(N4200), .C(N3913), .Y(N4447) );
  NAND2X1 gate1319_1 ( .A(N4305), .B(N4200), .Y(N4448_1) );
  NAND2X1 gate1319_2 ( .A(N4213), .B(N4167), .Y(N4448_2) );
  NAND2X1 gate1319 ( .A(N4448_1), .B(N4448_2), .Y(N4448) );
  INVX1 gate1320 ( .A(N4356), .Y(N4452) );
  NAND2X1 gate1321 ( .A(N4329), .B(N4393), .Y(N4458) );
  INVX1 gate1322 ( .A(N4365), .Y(N4461) );
  INVX1 gate1323 ( .A(N4368), .Y(N4462) );
  NAND2X1 gate1324 ( .A(N4371), .B(N1460), .Y(N4463) );
  INVX1 gate1325 ( .A(N4371), .Y(N4464) );
  BUFX2 gate1326 ( .A(N4310), .Y(N4465) );
  NOR2X1 gate1327 ( .A(N4331), .B(N4296), .Y(N4468) );
  AND2X1 gate1328 ( .A(N4376), .B(N2732), .Y(N4472) );
  AND2X1 gate1329 ( .A(N4377), .B(N2740), .Y(N4475) );
  BUFX2 gate1330 ( .A(N4310), .Y(N4479) );
  INVX1 gate1331 ( .A(N4353), .Y(N4484) );
  INVX1 gate1332 ( .A(N4359), .Y(N4486) );
  NAND2X1 gate1333 ( .A(N4359), .B(N4299), .Y(N4487) );
  INVX1 gate1334 ( .A(N4362), .Y(N4491) );
  AND2X1 gate1335 ( .A(N330), .B(N4319), .Y(N4493) );
  INVX1 gate1336 ( .A(N4398), .Y(N4496) );
  AND2X1 gate1337 ( .A(N4287), .B(N4398), .Y(N4497) );
  AND2X1 gate1338 ( .A(N4442), .B(N1769), .Y(N4498) );
  NAND2X1 gate1339_1 ( .A(N3947), .B(N4446), .Y(N4503_1) );
  NAND2X1 gate1339_2 ( .A(N4447), .B(N4448), .Y(N4503_2) );
  NAND2X1 gate1339 ( .A(N4503_1), .B(N4503_2), .Y(N4503) );
  INVX1 gate1340 ( .A(N4413), .Y(N4506) );
  INVX1 gate1341 ( .A(N4435), .Y(N4507) );
  INVX1 gate1342 ( .A(N4421), .Y(N4508) );
  NAND2X1 gate1343 ( .A(N4421), .B(N4452), .Y(N4509) );
  INVX1 gate1344 ( .A(N4427), .Y(N4510) );
  NAND2X1 gate1345 ( .A(N4427), .B(N4241), .Y(N4511) );
  NAND2X1 gate1346 ( .A(N965), .B(N4464), .Y(N4515) );
  INVX1 gate1347 ( .A(N4416), .Y(N4526) );
  NAND2X1 gate1348 ( .A(N4416), .B(N4484), .Y(N4527) );
  NAND2X1 gate1349 ( .A(N4182), .B(N4486), .Y(N4528) );
  INVX1 gate1350 ( .A(N4430), .Y(N4529) );
  NAND2X1 gate1351 ( .A(N4430), .B(N4491), .Y(N4530) );
  BUFX2 gate1352 ( .A(N4387), .Y(N4531) );
  BUFX2 gate1353 ( .A(N4387), .Y(N4534) );
  BUFX2 gate1354 ( .A(N4390), .Y(N4537) );
  BUFX2 gate1355 ( .A(N4390), .Y(N4540) );
  AND2X1 gate1356_1 ( .A(N330), .B(N4319), .Y(N4545_1) );
  AND2X1 gate1356 ( .A(N4496), .B(N4545_1), .Y(N4545) );
  AND2X1 gate1357 ( .A(N330), .B(N4443), .Y(N4549) );
  NAND2X1 gate1358 ( .A(N4356), .B(N4508), .Y(N4552) );
  NAND2X1 gate1359 ( .A(N4142), .B(N4510), .Y(N4555) );
  INVX1 gate1360 ( .A(N4493), .Y(N4558) );
  NAND2X1 gate1361 ( .A(N4463), .B(N4515), .Y(N4559) );
  INVX1 gate1362 ( .A(N4465), .Y(N4562) );
  AND2X1 gate1363 ( .A(N4310), .B(N4465), .Y(N4563) );
  BUFX2 gate1364 ( .A(N4468), .Y(N4564) );
  INVX1 gate1365 ( .A(N4479), .Y(N4568) );
  BUFX2 gate1366 ( .A(N4443), .Y(N4569) );
  NAND2X1 gate1367 ( .A(N4353), .B(N4526), .Y(N4572) );
  NAND2X1 gate1368 ( .A(N4362), .B(N4529), .Y(N4573) );
  NAND2X1 gate1369 ( .A(N4487), .B(N4528), .Y(N4576) );
  BUFX2 gate1370 ( .A(N4458), .Y(N4581) );
  BUFX2 gate1371 ( .A(N4458), .Y(N4584) );
  OR2X1 gate1372_1 ( .A(N2758), .B(N4498), .Y(N4587_1) );
  OR2X1 gate1372 ( .A(N2761), .B(N4587_1), .Y(N4587) );
  NOR3X1 gate1373 ( .A(N2758), .B(N4498), .C(N2761), .Y(N4588) );
  OR2X1 gate1374 ( .A(N4545), .B(N4497), .Y(N4589) );
  NAND2X1 gate1375 ( .A(N4552), .B(N4509), .Y(N4593) );
  INVX1 gate1376 ( .A(N4531), .Y(N4596) );
  INVX1 gate1377 ( .A(N4534), .Y(N4597) );
  NAND2X1 gate1378 ( .A(N4555), .B(N4511), .Y(N4599) );
  INVX1 gate1379 ( .A(N4537), .Y(N4602) );
  INVX1 gate1380 ( .A(N4540), .Y(N4603) );
  AND2X1 gate1381_1 ( .A(N330), .B(N4284), .Y(N4608_1) );
  AND2X1 gate1381 ( .A(N4562), .B(N4608_1), .Y(N4608) );
  BUFX2 gate1382 ( .A(N4503), .Y(N4613) );
  BUFX2 gate1383 ( .A(N4503), .Y(N4616) );
  NAND2X1 gate1384 ( .A(N4572), .B(N4527), .Y(N4619) );
  NAND2X1 gate1385 ( .A(N4573), .B(N4530), .Y(N4623) );
  INVX1 gate1386 ( .A(N4588), .Y(N4628) );
  NAND2X1 gate1387 ( .A(N4569), .B(N4506), .Y(N4629) );
  INVX1 gate1388 ( .A(N4569), .Y(N4630) );
  INVX1 gate1389 ( .A(N4576), .Y(N4635) );
  NAND2X1 gate1390 ( .A(N4576), .B(N4291), .Y(N4636) );
  INVX1 gate1391 ( .A(N4581), .Y(N4640) );
  NAND2X1 gate1392 ( .A(N4581), .B(N4461), .Y(N4641) );
  INVX1 gate1393 ( .A(N4584), .Y(N4642) );
  NAND2X1 gate1394 ( .A(N4584), .B(N4462), .Y(N4643) );
  NOR2X1 gate1395 ( .A(N4608), .B(N4563), .Y(N4644) );
  AND2X1 gate1396 ( .A(N4559), .B(N2128), .Y(N4647) );
  AND2X1 gate1397 ( .A(N4559), .B(N2743), .Y(N4650) );
  BUFX2 gate1398 ( .A(N4549), .Y(N4656) );
  BUFX2 gate1399 ( .A(N4549), .Y(N4659) );
  BUFX2 gate1400 ( .A(N4564), .Y(N4664) );
  AND2X1 gate1401 ( .A(N4587), .B(N4628), .Y(N4667) );
  NAND2X1 gate1402 ( .A(N4413), .B(N4630), .Y(N4668) );
  INVX1 gate1403 ( .A(N4616), .Y(N4669) );
  NAND2X1 gate1404 ( .A(N4616), .B(N4239), .Y(N4670) );
  INVX1 gate1405 ( .A(N4619), .Y(N4673) );
  NAND2X1 gate1406 ( .A(N4619), .B(N4507), .Y(N4674) );
  NAND2X1 gate1407 ( .A(N4186), .B(N4635), .Y(N4675) );
  INVX1 gate1408 ( .A(N4623), .Y(N4676) );
  NAND2X1 gate1409 ( .A(N4623), .B(N4558), .Y(N4677) );
  NAND2X1 gate1410 ( .A(N4365), .B(N4640), .Y(N4678) );
  NAND2X1 gate1411 ( .A(N4368), .B(N4642), .Y(N4679) );
  INVX1 gate1412 ( .A(N4613), .Y(N4687) );
  NAND2X1 gate1413 ( .A(N4613), .B(N4568), .Y(N4688) );
  BUFX2 gate1414 ( .A(N4593), .Y(N4691) );
  BUFX2 gate1415 ( .A(N4593), .Y(N4694) );
  BUFX2 gate1416 ( .A(N4599), .Y(N4697) );
  BUFX2 gate1417 ( .A(N4599), .Y(N4700) );
  NAND2X1 gate1418 ( .A(N4629), .B(N4668), .Y(N4704) );
  NAND2X1 gate1419 ( .A(N4139), .B(N4669), .Y(N4705) );
  INVX1 gate1420 ( .A(N4656), .Y(N4706) );
  INVX1 gate1421 ( .A(N4659), .Y(N4707) );
  NAND2X1 gate1422 ( .A(N4435), .B(N4673), .Y(N4708) );
  NAND2X1 gate1423 ( .A(N4675), .B(N4636), .Y(N4711) );
  NAND2X1 gate1424 ( .A(N4493), .B(N4676), .Y(N4716) );
  NAND2X1 gate1425 ( .A(N4678), .B(N4641), .Y(N4717) );
  NAND2X1 gate1426 ( .A(N4679), .B(N4643), .Y(N4721) );
  BUFX2 gate1427 ( .A(N4644), .Y(N4722) );
  INVX1 gate1428 ( .A(N4664), .Y(N4726) );
  OR2X1 gate1429_1 ( .A(N4647), .B(N4650), .Y(N4727_1) );
  OR2X1 gate1429 ( .A(N4350), .B(N4727_1), .Y(N4727) );
  NOR3X1 gate1430 ( .A(N4647), .B(N4650), .C(N4350), .Y(N4730) );
  NAND2X1 gate1431 ( .A(N4479), .B(N4687), .Y(N4733) );
  NAND2X1 gate1432 ( .A(N4705), .B(N4670), .Y(N4740) );
  NAND2X1 gate1433 ( .A(N4708), .B(N4674), .Y(N4743) );
  INVX1 gate1434 ( .A(N4691), .Y(N4747) );
  NAND2X1 gate1435 ( .A(N4691), .B(N4596), .Y(N4748) );
  INVX1 gate1436 ( .A(N4694), .Y(N4749) );
  NAND2X1 gate1437 ( .A(N4694), .B(N4597), .Y(N4750) );
  INVX1 gate1438 ( .A(N4697), .Y(N4753) );
  NAND2X1 gate1439 ( .A(N4697), .B(N4602), .Y(N4754) );
  INVX1 gate1440 ( .A(N4700), .Y(N4755) );
  NAND2X1 gate1441 ( .A(N4700), .B(N4603), .Y(N4756) );
  NAND2X1 gate1442 ( .A(N4716), .B(N4677), .Y(N4757) );
  NAND2X1 gate1443 ( .A(N4733), .B(N4688), .Y(N4769) );
  AND2X1 gate1444 ( .A(N330), .B(N4704), .Y(N4772) );
  INVX1 gate1445 ( .A(N4721), .Y(N4775) );
  INVX1 gate1446 ( .A(N4730), .Y(N4778) );
  NAND2X1 gate1447 ( .A(N4531), .B(N4747), .Y(N4786) );
  NAND2X1 gate1448 ( .A(N4534), .B(N4749), .Y(N4787) );
  NAND2X1 gate1449 ( .A(N4537), .B(N4753), .Y(N4788) );
  NAND2X1 gate1450 ( .A(N4540), .B(N4755), .Y(N4789) );
  AND2X1 gate1451 ( .A(N4711), .B(N2124), .Y(N4794) );
  AND2X1 gate1452 ( .A(N4711), .B(N2735), .Y(N4797) );
  AND2X1 gate1453 ( .A(N4717), .B(N2127), .Y(N4800) );
  BUFX2 gate1454 ( .A(N4722), .Y(N4805) );
  AND2X1 gate1455 ( .A(N4717), .B(N4468), .Y(N4808) );
  BUFX2 gate1456 ( .A(N4727), .Y(N4812) );
  AND2X1 gate1457 ( .A(N4727), .B(N4778), .Y(N4815) );
  INVX1 gate1458 ( .A(N4769), .Y(N4816) );
  INVX1 gate1459 ( .A(N4772), .Y(N4817) );
  NAND2X1 gate1460 ( .A(N4786), .B(N4748), .Y(N4818) );
  NAND2X1 gate1461 ( .A(N4787), .B(N4750), .Y(N4822) );
  NAND2X1 gate1462 ( .A(N4788), .B(N4754), .Y(N4823) );
  NAND2X1 gate1463 ( .A(N4789), .B(N4756), .Y(N4826) );
  NAND2X1 gate1464 ( .A(N4775), .B(N4726), .Y(N4829) );
  INVX1 gate1465 ( .A(N4775), .Y(N4830) );
  AND2X1 gate1466 ( .A(N4743), .B(N2122), .Y(N4831) );
  AND2X1 gate1467 ( .A(N4757), .B(N2126), .Y(N4838) );
  BUFX2 gate1468 ( .A(N4740), .Y(N4844) );
  BUFX2 gate1469 ( .A(N4740), .Y(N4847) );
  BUFX2 gate1470 ( .A(N4743), .Y(N4850) );
  BUFX2 gate1471 ( .A(N4757), .Y(N4854) );
  NAND2X1 gate1472 ( .A(N4772), .B(N4816), .Y(N4859) );
  NAND2X1 gate1473 ( .A(N4769), .B(N4817), .Y(N4860) );
  INVX1 gate1474 ( .A(N4826), .Y(N4868) );
  INVX1 gate1475 ( .A(N4805), .Y(N4870) );
  INVX1 gate1476 ( .A(N4808), .Y(N4872) );
  NAND2X1 gate1477 ( .A(N4664), .B(N4830), .Y(N4873) );
  OR2X1 gate1478_1 ( .A(N4794), .B(N4797), .Y(N4876_1) );
  OR2X1 gate1478 ( .A(N4341), .B(N4876_1), .Y(N4876) );
  NOR3X1 gate1479 ( .A(N4794), .B(N4797), .C(N4341), .Y(N4880) );
  INVX1 gate1480 ( .A(N4812), .Y(N4885) );
  INVX1 gate1481 ( .A(N4822), .Y(N4889) );
  NAND2X1 gate1482 ( .A(N4859), .B(N4860), .Y(N4895) );
  INVX1 gate1483 ( .A(N4844), .Y(N4896) );
  NAND2X1 gate1484 ( .A(N4844), .B(N4706), .Y(N4897) );
  INVX1 gate1485 ( .A(N4847), .Y(N4898) );
  NAND2X1 gate1486 ( .A(N4847), .B(N4707), .Y(N4899) );
  NOR2X1 gate1487 ( .A(N4868), .B(N4564), .Y(N4900) );
  AND2X1 gate1488_1 ( .A(N4717), .B(N4757), .Y(N4901_1) );
  AND2X1 gate1488_2 ( .A(N4823), .B(N4564), .Y(N4901_2) );
  AND2X1 gate1488 ( .A(N4901_1), .B(N4901_2), .Y(N4901) );
  INVX1 gate1489 ( .A(N4850), .Y(N4902) );
  INVX1 gate1490 ( .A(N4854), .Y(N4904) );
  NAND2X1 gate1491 ( .A(N4854), .B(N4872), .Y(N4905) );
  NAND2X1 gate1492 ( .A(N4873), .B(N4829), .Y(N4906) );
  AND2X1 gate1493 ( .A(N4818), .B(N2123), .Y(N4907) );
  AND2X1 gate1494 ( .A(N4823), .B(N2125), .Y(N4913) );
  AND2X1 gate1495 ( .A(N4818), .B(N4644), .Y(N4916) );
  INVX1 gate1496 ( .A(N4880), .Y(N4920) );
  AND2X1 gate1497 ( .A(N4895), .B(N2184), .Y(N4921) );
  NAND2X1 gate1498 ( .A(N4656), .B(N4896), .Y(N4924) );
  NAND2X1 gate1499 ( .A(N4659), .B(N4898), .Y(N4925) );
  OR2X1 gate1500 ( .A(N4900), .B(N4901), .Y(N4926) );
  NAND2X1 gate1501 ( .A(N4889), .B(N4870), .Y(N4928) );
  INVX1 gate1502 ( .A(N4889), .Y(N4929) );
  NAND2X1 gate1503 ( .A(N4808), .B(N4904), .Y(N4930) );
  INVX1 gate1504 ( .A(N4906), .Y(N4931) );
  BUFX2 gate1505 ( .A(N4876), .Y(N4937) );
  BUFX2 gate1506 ( .A(N4876), .Y(N4940) );
  AND2X1 gate1507 ( .A(N4876), .B(N4920), .Y(N4944) );
  NAND2X1 gate1508 ( .A(N4924), .B(N4897), .Y(N4946) );
  NAND2X1 gate1509 ( .A(N4925), .B(N4899), .Y(N4949) );
  NAND2X1 gate1510 ( .A(N4916), .B(N4902), .Y(N4950) );
  INVX1 gate1511 ( .A(N4916), .Y(N4951) );
  NAND2X1 gate1512 ( .A(N4805), .B(N4929), .Y(N4952) );
  NAND2X1 gate1513 ( .A(N4930), .B(N4905), .Y(N4953) );
  AND2X1 gate1514 ( .A(N4926), .B(N2737), .Y(N4954) );
  AND2X1 gate1515 ( .A(N4931), .B(N2741), .Y(N4957) );
  OR2X1 gate1516_1 ( .A(N2764), .B(N2483), .Y(N4964_1) );
  OR2X1 gate1516 ( .A(N4921), .B(N4964_1), .Y(N4964) );
  NOR3X1 gate1517 ( .A(N2764), .B(N2483), .C(N4921), .Y(N4965) );
  INVX1 gate1518 ( .A(N4949), .Y(N4968) );
  NAND2X1 gate1519 ( .A(N4850), .B(N4951), .Y(N4969) );
  NAND2X1 gate1520 ( .A(N4952), .B(N4928), .Y(N4970) );
  AND2X1 gate1521 ( .A(N4953), .B(N2739), .Y(N4973) );
  INVX1 gate1522 ( .A(N4937), .Y(N4978) );
  INVX1 gate1523 ( .A(N4940), .Y(N4979) );
  INVX1 gate1524 ( .A(N4965), .Y(N4980) );
  NOR2X1 gate1525 ( .A(N4968), .B(N4722), .Y(N4981) );
  AND2X1 gate1526_1 ( .A(N4818), .B(N4743), .Y(N4982_1) );
  AND2X1 gate1526_2 ( .A(N4946), .B(N4722), .Y(N4982_2) );
  AND2X1 gate1526 ( .A(N4982_1), .B(N4982_2), .Y(N4982) );
  NAND2X1 gate1527 ( .A(N4950), .B(N4969), .Y(N4983) );
  INVX1 gate1528 ( .A(N4970), .Y(N4984) );
  AND2X1 gate1529 ( .A(N4946), .B(N2121), .Y(N4985) );
  OR2X1 gate1530_1 ( .A(N4913), .B(N4954), .Y(N4988_1) );
  OR2X1 gate1530 ( .A(N4344), .B(N4988_1), .Y(N4988) );
  NOR3X1 gate1531 ( .A(N4913), .B(N4954), .C(N4344), .Y(N4991) );
  OR2X1 gate1532_1 ( .A(N4800), .B(N4957), .Y(N4996_1) );
  OR2X1 gate1532 ( .A(N4347), .B(N4996_1), .Y(N4996) );
  NOR3X1 gate1533 ( .A(N4800), .B(N4957), .C(N4347), .Y(N4999) );
  AND2X1 gate1534 ( .A(N4964), .B(N4980), .Y(N5002) );
  OR2X1 gate1535 ( .A(N4981), .B(N4982), .Y(N5007) );
  AND2X1 gate1536 ( .A(N4983), .B(N2731), .Y(N5010) );
  AND2X1 gate1537 ( .A(N4984), .B(N2733), .Y(N5013) );
  OR2X1 gate1538_1 ( .A(N4838), .B(N4973), .Y(N5018_1) );
  OR2X1 gate1538 ( .A(N4475), .B(N5018_1), .Y(N5018) );
  NOR3X1 gate1539 ( .A(N4838), .B(N4973), .C(N4475), .Y(N5021) );
  INVX1 gate1540 ( .A(N4991), .Y(N5026) );
  INVX1 gate1541 ( .A(N4999), .Y(N5029) );
  AND2X1 gate1542 ( .A(N5007), .B(N2729), .Y(N5030) );
  BUFX2 gate1543 ( .A(N4996), .Y(N5039) );
  BUFX2 gate1544 ( .A(N4988), .Y(N5042) );
  AND2X1 gate1545 ( .A(N4988), .B(N5026), .Y(N5045) );
  INVX1 gate1546 ( .A(N5021), .Y(N5046) );
  AND2X1 gate1547 ( .A(N4996), .B(N5029), .Y(N5047) );
  OR2X1 gate1548_1 ( .A(N4831), .B(N5010), .Y(N5050_1) );
  OR2X1 gate1548 ( .A(N4472), .B(N5050_1), .Y(N5050) );
  NOR3X1 gate1549 ( .A(N4831), .B(N5010), .C(N4472), .Y(N5055) );
  OR2X1 gate1550_1 ( .A(N4907), .B(N5013), .Y(N5058_1) );
  OR2X1 gate1550 ( .A(N4338), .B(N5058_1), .Y(N5058) );
  NOR3X1 gate1551 ( .A(N4907), .B(N5013), .C(N4338), .Y(N5061) );
  AND2X1 gate1552_1 ( .A(N4730), .B(N4999), .Y(N5066_1) );
  AND2X1 gate1552_2 ( .A(N5021), .B(N4991), .Y(N5066_2) );
  AND2X1 gate1552 ( .A(N5066_1), .B(N5066_2), .Y(N5066) );
  BUFX2 gate1553 ( .A(N5018), .Y(N5070) );
  AND2X1 gate1554 ( .A(N5018), .B(N5046), .Y(N5078) );
  OR2X1 gate1555_1 ( .A(N4985), .B(N5030), .Y(N5080_1) );
  OR2X1 gate1555 ( .A(N4335), .B(N5080_1), .Y(N5080) );
  NOR3X1 gate1556 ( .A(N4985), .B(N5030), .C(N4335), .Y(N5085) );
  NAND2X1 gate1557 ( .A(N5039), .B(N4885), .Y(N5094) );
  INVX1 gate1558 ( .A(N5039), .Y(N5095) );
  INVX1 gate1559 ( .A(N5042), .Y(N5097) );
  AND2X1 gate1560 ( .A(N5050), .B(N5050), .Y(N5102) );
  INVX1 gate1561 ( .A(N5061), .Y(N5103) );
  NAND2X1 gate1562 ( .A(N4812), .B(N5095), .Y(N5108) );
  INVX1 gate1563 ( .A(N5070), .Y(N5109) );
  NAND2X1 gate1564 ( .A(N5070), .B(N5097), .Y(N5110) );
  BUFX2 gate1565 ( .A(N5058), .Y(N5111) );
  AND2X1 gate1566 ( .A(N5050), .B(N1461), .Y(N5114) );
  BUFX2 gate1567 ( .A(N5050), .Y(N5117) );
  AND2X1 gate1568 ( .A(N5080), .B(N5080), .Y(N5120) );
  AND2X1 gate1569 ( .A(N5058), .B(N5103), .Y(N5121) );
  NAND2X1 gate1570 ( .A(N5094), .B(N5108), .Y(N5122) );
  NAND2X1 gate1571 ( .A(N5042), .B(N5109), .Y(N5125) );
  AND2X1 gate1572 ( .A(N1461), .B(N5080), .Y(N5128) );
  AND2X1 gate1573_1 ( .A(N4880), .B(N5061), .Y(N5133_1) );
  AND2X1 gate1573_2 ( .A(N5055), .B(N5085), .Y(N5133_2) );
  AND2X1 gate1573 ( .A(N5133_1), .B(N5133_2), .Y(N5133) );
  AND2X1 gate1574_1 ( .A(N5055), .B(N5085), .Y(N5136_1) );
  AND2X1 gate1574 ( .A(N1464), .B(N5136_1), .Y(N5136) );
  BUFX2 gate1575 ( .A(N5080), .Y(N5139) );
  NAND2X1 gate1576 ( .A(N5125), .B(N5110), .Y(N5145) );
  BUFX2 gate1577 ( .A(N5111), .Y(N5151) );
  BUFX2 gate1578 ( .A(N5111), .Y(N5154) );
  INVX1 gate1579 ( .A(N5117), .Y(N5159) );
  BUFX2 gate1580 ( .A(N5114), .Y(N5160) );
  BUFX2 gate1581 ( .A(N5114), .Y(N5163) );
  AND2X1 gate1582 ( .A(N5066), .B(N5133), .Y(N5166) );
  AND2X1 gate1583 ( .A(N5066), .B(N5133), .Y(N5173) );
  BUFX2 gate1584 ( .A(N5122), .Y(N5174) );
  BUFX2 gate1585 ( .A(N5122), .Y(N5177) );
  INVX1 gate1586 ( .A(N5139), .Y(N5182) );
  NAND2X1 gate1587 ( .A(N5139), .B(N5159), .Y(N5183) );
  BUFX2 gate1588 ( .A(N5128), .Y(N5184) );
  BUFX2 gate1589 ( .A(N5128), .Y(N5188) );
  INVX1 gate1590 ( .A(N5166), .Y(N5192) );
  NOR2X1 gate1591 ( .A(N5136), .B(N5173), .Y(N5193) );
  NAND2X1 gate1592 ( .A(N5151), .B(N4978), .Y(N5196) );
  INVX1 gate1593 ( .A(N5151), .Y(N5197) );
  NAND2X1 gate1594 ( .A(N5154), .B(N4979), .Y(N5198) );
  INVX1 gate1595 ( .A(N5154), .Y(N5199) );
  INVX1 gate1596 ( .A(N5160), .Y(N5201) );
  INVX1 gate1597 ( .A(N5163), .Y(N5203) );
  BUFX2 gate1598 ( .A(N5145), .Y(N5205) );
  BUFX2 gate1599 ( .A(N5145), .Y(N5209) );
  NAND2X1 gate1600 ( .A(N5117), .B(N5182), .Y(N5212) );
  AND2X1 gate1601 ( .A(N213), .B(N5193), .Y(N5215) );
  INVX1 gate1602 ( .A(N5174), .Y(N5217) );
  INVX1 gate1603 ( .A(N5177), .Y(N5219) );
  NAND2X1 gate1604 ( .A(N4937), .B(N5197), .Y(N5220) );
  NAND2X1 gate1605 ( .A(N4940), .B(N5199), .Y(N5221) );
  INVX1 gate1606 ( .A(N5184), .Y(N5222) );
  NAND2X1 gate1607 ( .A(N5184), .B(N5201), .Y(N5223) );
  NAND2X1 gate1608 ( .A(N5188), .B(N5203), .Y(N5224) );
  INVX1 gate1609 ( .A(N5188), .Y(N5225) );
  NAND2X1 gate1610 ( .A(N5183), .B(N5212), .Y(N5228) );
  INVX1 gate1611 ( .A(N5215), .Y(N5231) );
  NAND2X1 gate1612 ( .A(N5205), .B(N5217), .Y(N5232) );
  INVX1 gate1613 ( .A(N5205), .Y(N5233) );
  NAND2X1 gate1614 ( .A(N5209), .B(N5219), .Y(N5234) );
  INVX1 gate1615 ( .A(N5209), .Y(N5235) );
  NAND2X1 gate1616 ( .A(N5196), .B(N5220), .Y(N5236) );
  NAND2X1 gate1617 ( .A(N5198), .B(N5221), .Y(N5240) );
  NAND2X1 gate1618 ( .A(N5160), .B(N5222), .Y(N5242) );
  NAND2X1 gate1619 ( .A(N5163), .B(N5225), .Y(N5243) );
  NAND2X1 gate1620 ( .A(N5174), .B(N5233), .Y(N5245) );
  NAND2X1 gate1621 ( .A(N5177), .B(N5235), .Y(N5246) );
  INVX1 gate1622 ( .A(N5240), .Y(N5250) );
  INVX1 gate1623 ( .A(N5228), .Y(N5253) );
  NAND2X1 gate1624 ( .A(N5242), .B(N5223), .Y(N5254) );
  NAND2X1 gate1625 ( .A(N5243), .B(N5224), .Y(N5257) );
  NAND2X1 gate1626 ( .A(N5232), .B(N5245), .Y(N5258) );
  NAND2X1 gate1627 ( .A(N5234), .B(N5246), .Y(N5261) );
  INVX1 gate1628 ( .A(N5257), .Y(N5266) );
  BUFX2 gate1629 ( .A(N5236), .Y(N5269) );
  AND2X1 gate1630_1 ( .A(N5236), .B(N5254), .Y(N5277_1) );
  AND2X1 gate1630 ( .A(N2307), .B(N5277_1), .Y(N5277) );
  AND2X1 gate1631_1 ( .A(N5250), .B(N5254), .Y(N5278_1) );
  AND2X1 gate1631 ( .A(N2310), .B(N5278_1), .Y(N5278) );
  INVX1 gate1632 ( .A(N5261), .Y(N5279) );
  INVX1 gate1633 ( .A(N5269), .Y(N5283) );
  NAND2X1 gate1634 ( .A(N5269), .B(N5253), .Y(N5284) );
  AND2X1 gate1635_1 ( .A(N5236), .B(N5266), .Y(N5285_1) );
  AND2X1 gate1635 ( .A(N2310), .B(N5285_1), .Y(N5285) );
  AND2X1 gate1636_1 ( .A(N5250), .B(N5266), .Y(N5286_1) );
  AND2X1 gate1636 ( .A(N2307), .B(N5286_1), .Y(N5286) );
  BUFX2 gate1637 ( .A(N5258), .Y(N5289) );
  BUFX2 gate1638 ( .A(N5258), .Y(N5292) );
  NAND2X1 gate1639 ( .A(N5228), .B(N5283), .Y(N5295) );
  OR2X1 gate1640_1 ( .A(N5277), .B(N5285), .Y(N5298_1) );
  OR2X1 gate1640_2 ( .A(N5278), .B(N5286), .Y(N5298_2) );
  OR2X1 gate1640 ( .A(N5298_1), .B(N5298_2), .Y(N5298) );
  BUFX2 gate1641 ( .A(N5279), .Y(N5303) );
  BUFX2 gate1642 ( .A(N5279), .Y(N5306) );
  NAND2X1 gate1643 ( .A(N5295), .B(N5284), .Y(N5309) );
  INVX1 gate1644 ( .A(N5292), .Y(N5312) );
  INVX1 gate1645 ( .A(N5289), .Y(N5313) );
  INVX1 gate1646 ( .A(N5306), .Y(N5322) );
  INVX1 gate1647 ( .A(N5303), .Y(N5323) );
  BUFX2 gate1648 ( .A(N5298), .Y(N5324) );
  BUFX2 gate1649 ( .A(N5298), .Y(N5327) );
  BUFX2 gate1650 ( .A(N5309), .Y(N5332) );
  BUFX2 gate1651 ( .A(N5309), .Y(N5335) );
  NAND2X1 gate1652 ( .A(N5324), .B(N5323), .Y(N5340) );
  NAND2X1 gate1653 ( .A(N5327), .B(N5322), .Y(N5341) );
  INVX1 gate1654 ( .A(N5327), .Y(N5344) );
  INVX1 gate1655 ( .A(N5324), .Y(N5345) );
  NAND2X1 gate1656 ( .A(N5332), .B(N5313), .Y(N5348) );
  NAND2X1 gate1657 ( .A(N5335), .B(N5312), .Y(N5349) );
  NAND2X1 gate1658 ( .A(N5303), .B(N5345), .Y(N5350) );
  NAND2X1 gate1659 ( .A(N5306), .B(N5344), .Y(N5351) );
  INVX1 gate1660 ( .A(N5335), .Y(N5352) );
  INVX1 gate1661 ( .A(N5332), .Y(N5353) );
  NAND2X1 gate1662 ( .A(N5289), .B(N5353), .Y(N5354) );
  NAND2X1 gate1663 ( .A(N5292), .B(N5352), .Y(N5355) );
  NAND2X1 gate1664 ( .A(N5350), .B(N5340), .Y(N5356) );
  NAND2X1 gate1665 ( .A(N5351), .B(N5341), .Y(N5357) );
  NAND2X1 gate1666 ( .A(N5348), .B(N5354), .Y(N5358) );
  NAND2X1 gate1667 ( .A(N5349), .B(N5355), .Y(N5359) );
  AND2X1 gate1668 ( .A(N5356), .B(N5357), .Y(N5360) );
  NAND2X1 gate1669 ( .A(N5358), .B(N5359), .Y(N5361) );
endmodule



module c1355_synth ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272,
         G275, G278, G281, G284, G287, G290, G293, G296, G299, G302, G305,
         G308, G311, G314, G317, G320, G323, G326, G329, G332, G335, G338,
         G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365,
         G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376,
         G377, G378, G379, G380, G381, G382, G383, G384, G385, G386, G387,
         G388, G389, G390, G391, G392, G393, G394, G395, G396, G397, G398,
         G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409,
         G410, G411, G412, G413, G414, G415, G416, G417, G418, G419, G420,
         G421, G422, G423, G424, G425, G426, G429, G432, G435, G438, G441,
         G444, G447, G450, G453, G456, G459, G462, G465, G468, G471, G474,
         G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507,
         G510, G513, G516, G519, G522, G525, G528, G531, G534, G537, G540,
         G543, G546, G549, G552, G555, G558, G561, G564, G567, G570, G571,
         G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, G582,
         G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593,
         G594, G595, G596, G597, G598, G599, G600, G601, G602, G607, G612,
         G617, G622, G627, G632, G637, G642, G645, G648, G651, G654, G657,
         G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690,
         G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701,
         G702, G703, G704, G705, G706, G709, G712, G715, G718, G721, G724,
         G727, G730, G733, G736, G739, G742, G745, G748, G751, G754, G755,
         G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766,
         G767, G768, G769, G770, G773, G776, G779, G782, G785, G788, G791,
         G794, G797, G800, G803, G806, G809, G812, G815, G818, G819, G820,
         G821, G822, G823, G824, G825, G826, G827, G828, G829, G830, G831,
         G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938,
         G939, G940, G941, G942, G943, G944, G945, G946, G947, G948, G949,
         G950, G951, G952, G953, G954, G955, G956, G957, G958, G959, G960,
         G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, G971,
         G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982,
         G983, G984, G985, G986, G991, G996, G1001, G1006, G1011, G1016, G1021,
         G1026, G1031, G1036, G1039, G1042, G1045, G1048, G1051, G1054, G1057,
         G1060, G1063, G1066, G1069, G1072, G1075, G1078, G1081, G1084, G1087,
         G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, G1117,
         G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147,
         G1150, G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177,
         G1180, G1183, G1186, G1189, G1192, G1195, G1198, G1201, G1204, G1207,
         G1210, G1213, G1216, G1219, G1222, G1225, G1228, G1229, G1230, G1231,
         G1232, G1233, G1234, G1235, G1236, G1237, G1238, G1239, G1240, G1241,
         G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, G1251,
         G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261,
         G1262, G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271,
         G1272, G1273, G1274, G1275, G1276, G1277, G1278, G1279, G1280, G1281,
         G1282, G1283, G1284, G1285, G1286, G1287, G1288, G1289, G1290, G1291,
         G1292, G1293, G1294, G1295, G1296, G1297, G1298, G1299, G1300, G1301,
         G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, G1311,
         G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321,
         G1322, G1323, G978_1, G978_2, G979_1, G979_2, G980_1, G980_2, G981_1,
         G981_2, G982_1, G982_2, G983_1, G983_2, G984_1, G984_2, G985_1,
         G985_2, G986_1, G986_2, G991_1, G991_2, G996_1, G996_2, G996_3,
         G1001_1, G1001_2, G1001_3, G1006_1, G1006_2, G1006_3, G1011_1,
         G1011_2, G1011_3, G1016_1, G1016_2, G1016_3, G1021_1, G1021_2,
         G1021_3, G1026_1, G1026_2, G1026_3, G1031_1, G1031_2, G1031_3;

  AND2X1 gate1 ( .A(G33), .B(G41), .Y(G242) );
  AND2X1 gate2 ( .A(G34), .B(G41), .Y(G245) );
  AND2X1 gate3 ( .A(G35), .B(G41), .Y(G248) );
  AND2X1 gate4 ( .A(G36), .B(G41), .Y(G251) );
  AND2X1 gate5 ( .A(G37), .B(G41), .Y(G254) );
  AND2X1 gate6 ( .A(G38), .B(G41), .Y(G257) );
  AND2X1 gate7 ( .A(G39), .B(G41), .Y(G260) );
  AND2X1 gate8 ( .A(G40), .B(G41), .Y(G263) );
  NAND2X1 gate9 ( .A(G1), .B(G2), .Y(G266) );
  NAND2X1 gate10 ( .A(G3), .B(G4), .Y(G269) );
  NAND2X1 gate11 ( .A(G5), .B(G6), .Y(G272) );
  NAND2X1 gate12 ( .A(G7), .B(G8), .Y(G275) );
  NAND2X1 gate13 ( .A(G9), .B(G10), .Y(G278) );
  NAND2X1 gate14 ( .A(G11), .B(G12), .Y(G281) );
  NAND2X1 gate15 ( .A(G13), .B(G14), .Y(G284) );
  NAND2X1 gate16 ( .A(G15), .B(G16), .Y(G287) );
  NAND2X1 gate17 ( .A(G17), .B(G18), .Y(G290) );
  NAND2X1 gate18 ( .A(G19), .B(G20), .Y(G293) );
  NAND2X1 gate19 ( .A(G21), .B(G22), .Y(G296) );
  NAND2X1 gate20 ( .A(G23), .B(G24), .Y(G299) );
  NAND2X1 gate21 ( .A(G25), .B(G26), .Y(G302) );
  NAND2X1 gate22 ( .A(G27), .B(G28), .Y(G305) );
  NAND2X1 gate23 ( .A(G29), .B(G30), .Y(G308) );
  NAND2X1 gate24 ( .A(G31), .B(G32), .Y(G311) );
  NAND2X1 gate25 ( .A(G1), .B(G5), .Y(G314) );
  NAND2X1 gate26 ( .A(G9), .B(G13), .Y(G317) );
  NAND2X1 gate27 ( .A(G2), .B(G6), .Y(G320) );
  NAND2X1 gate28 ( .A(G10), .B(G14), .Y(G323) );
  NAND2X1 gate29 ( .A(G3), .B(G7), .Y(G326) );
  NAND2X1 gate30 ( .A(G11), .B(G15), .Y(G329) );
  NAND2X1 gate31 ( .A(G4), .B(G8), .Y(G332) );
  NAND2X1 gate32 ( .A(G12), .B(G16), .Y(G335) );
  NAND2X1 gate33 ( .A(G17), .B(G21), .Y(G338) );
  NAND2X1 gate34 ( .A(G25), .B(G29), .Y(G341) );
  NAND2X1 gate35 ( .A(G18), .B(G22), .Y(G344) );
  NAND2X1 gate36 ( .A(G26), .B(G30), .Y(G347) );
  NAND2X1 gate37 ( .A(G19), .B(G23), .Y(G350) );
  NAND2X1 gate38 ( .A(G27), .B(G31), .Y(G353) );
  NAND2X1 gate39 ( .A(G20), .B(G24), .Y(G356) );
  NAND2X1 gate40 ( .A(G28), .B(G32), .Y(G359) );
  NAND2X1 gate41 ( .A(G1), .B(G266), .Y(G362) );
  NAND2X1 gate42 ( .A(G2), .B(G266), .Y(G363) );
  NAND2X1 gate43 ( .A(G3), .B(G269), .Y(G364) );
  NAND2X1 gate44 ( .A(G4), .B(G269), .Y(G365) );
  NAND2X1 gate45 ( .A(G5), .B(G272), .Y(G366) );
  NAND2X1 gate46 ( .A(G6), .B(G272), .Y(G367) );
  NAND2X1 gate47 ( .A(G7), .B(G275), .Y(G368) );
  NAND2X1 gate48 ( .A(G8), .B(G275), .Y(G369) );
  NAND2X1 gate49 ( .A(G9), .B(G278), .Y(G370) );
  NAND2X1 gate50 ( .A(G10), .B(G278), .Y(G371) );
  NAND2X1 gate51 ( .A(G11), .B(G281), .Y(G372) );
  NAND2X1 gate52 ( .A(G12), .B(G281), .Y(G373) );
  NAND2X1 gate53 ( .A(G13), .B(G284), .Y(G374) );
  NAND2X1 gate54 ( .A(G14), .B(G284), .Y(G375) );
  NAND2X1 gate55 ( .A(G15), .B(G287), .Y(G376) );
  NAND2X1 gate56 ( .A(G16), .B(G287), .Y(G377) );
  NAND2X1 gate57 ( .A(G17), .B(G290), .Y(G378) );
  NAND2X1 gate58 ( .A(G18), .B(G290), .Y(G379) );
  NAND2X1 gate59 ( .A(G19), .B(G293), .Y(G380) );
  NAND2X1 gate60 ( .A(G20), .B(G293), .Y(G381) );
  NAND2X1 gate61 ( .A(G21), .B(G296), .Y(G382) );
  NAND2X1 gate62 ( .A(G22), .B(G296), .Y(G383) );
  NAND2X1 gate63 ( .A(G23), .B(G299), .Y(G384) );
  NAND2X1 gate64 ( .A(G24), .B(G299), .Y(G385) );
  NAND2X1 gate65 ( .A(G25), .B(G302), .Y(G386) );
  NAND2X1 gate66 ( .A(G26), .B(G302), .Y(G387) );
  NAND2X1 gate67 ( .A(G27), .B(G305), .Y(G388) );
  NAND2X1 gate68 ( .A(G28), .B(G305), .Y(G389) );
  NAND2X1 gate69 ( .A(G29), .B(G308), .Y(G390) );
  NAND2X1 gate70 ( .A(G30), .B(G308), .Y(G391) );
  NAND2X1 gate71 ( .A(G31), .B(G311), .Y(G392) );
  NAND2X1 gate72 ( .A(G32), .B(G311), .Y(G393) );
  NAND2X1 gate73 ( .A(G1), .B(G314), .Y(G394) );
  NAND2X1 gate74 ( .A(G5), .B(G314), .Y(G395) );
  NAND2X1 gate75 ( .A(G9), .B(G317), .Y(G396) );
  NAND2X1 gate76 ( .A(G13), .B(G317), .Y(G397) );
  NAND2X1 gate77 ( .A(G2), .B(G320), .Y(G398) );
  NAND2X1 gate78 ( .A(G6), .B(G320), .Y(G399) );
  NAND2X1 gate79 ( .A(G10), .B(G323), .Y(G400) );
  NAND2X1 gate80 ( .A(G14), .B(G323), .Y(G401) );
  NAND2X1 gate81 ( .A(G3), .B(G326), .Y(G402) );
  NAND2X1 gate82 ( .A(G7), .B(G326), .Y(G403) );
  NAND2X1 gate83 ( .A(G11), .B(G329), .Y(G404) );
  NAND2X1 gate84 ( .A(G15), .B(G329), .Y(G405) );
  NAND2X1 gate85 ( .A(G4), .B(G332), .Y(G406) );
  NAND2X1 gate86 ( .A(G8), .B(G332), .Y(G407) );
  NAND2X1 gate87 ( .A(G12), .B(G335), .Y(G408) );
  NAND2X1 gate88 ( .A(G16), .B(G335), .Y(G409) );
  NAND2X1 gate89 ( .A(G17), .B(G338), .Y(G410) );
  NAND2X1 gate90 ( .A(G21), .B(G338), .Y(G411) );
  NAND2X1 gate91 ( .A(G25), .B(G341), .Y(G412) );
  NAND2X1 gate92 ( .A(G29), .B(G341), .Y(G413) );
  NAND2X1 gate93 ( .A(G18), .B(G344), .Y(G414) );
  NAND2X1 gate94 ( .A(G22), .B(G344), .Y(G415) );
  NAND2X1 gate95 ( .A(G26), .B(G347), .Y(G416) );
  NAND2X1 gate96 ( .A(G30), .B(G347), .Y(G417) );
  NAND2X1 gate97 ( .A(G19), .B(G350), .Y(G418) );
  NAND2X1 gate98 ( .A(G23), .B(G350), .Y(G419) );
  NAND2X1 gate99 ( .A(G27), .B(G353), .Y(G420) );
  NAND2X1 gate100 ( .A(G31), .B(G353), .Y(G421) );
  NAND2X1 gate101 ( .A(G20), .B(G356), .Y(G422) );
  NAND2X1 gate102 ( .A(G24), .B(G356), .Y(G423) );
  NAND2X1 gate103 ( .A(G28), .B(G359), .Y(G424) );
  NAND2X1 gate104 ( .A(G32), .B(G359), .Y(G425) );
  NAND2X1 gate105 ( .A(G362), .B(G363), .Y(G426) );
  NAND2X1 gate106 ( .A(G364), .B(G365), .Y(G429) );
  NAND2X1 gate107 ( .A(G366), .B(G367), .Y(G432) );
  NAND2X1 gate108 ( .A(G368), .B(G369), .Y(G435) );
  NAND2X1 gate109 ( .A(G370), .B(G371), .Y(G438) );
  NAND2X1 gate110 ( .A(G372), .B(G373), .Y(G441) );
  NAND2X1 gate111 ( .A(G374), .B(G375), .Y(G444) );
  NAND2X1 gate112 ( .A(G376), .B(G377), .Y(G447) );
  NAND2X1 gate113 ( .A(G378), .B(G379), .Y(G450) );
  NAND2X1 gate114 ( .A(G380), .B(G381), .Y(G453) );
  NAND2X1 gate115 ( .A(G382), .B(G383), .Y(G456) );
  NAND2X1 gate116 ( .A(G384), .B(G385), .Y(G459) );
  NAND2X1 gate117 ( .A(G386), .B(G387), .Y(G462) );
  NAND2X1 gate118 ( .A(G388), .B(G389), .Y(G465) );
  NAND2X1 gate119 ( .A(G390), .B(G391), .Y(G468) );
  NAND2X1 gate120 ( .A(G392), .B(G393), .Y(G471) );
  NAND2X1 gate121 ( .A(G394), .B(G395), .Y(G474) );
  NAND2X1 gate122 ( .A(G396), .B(G397), .Y(G477) );
  NAND2X1 gate123 ( .A(G398), .B(G399), .Y(G480) );
  NAND2X1 gate124 ( .A(G400), .B(G401), .Y(G483) );
  NAND2X1 gate125 ( .A(G402), .B(G403), .Y(G486) );
  NAND2X1 gate126 ( .A(G404), .B(G405), .Y(G489) );
  NAND2X1 gate127 ( .A(G406), .B(G407), .Y(G492) );
  NAND2X1 gate128 ( .A(G408), .B(G409), .Y(G495) );
  NAND2X1 gate129 ( .A(G410), .B(G411), .Y(G498) );
  NAND2X1 gate130 ( .A(G412), .B(G413), .Y(G501) );
  NAND2X1 gate131 ( .A(G414), .B(G415), .Y(G504) );
  NAND2X1 gate132 ( .A(G416), .B(G417), .Y(G507) );
  NAND2X1 gate133 ( .A(G418), .B(G419), .Y(G510) );
  NAND2X1 gate134 ( .A(G420), .B(G421), .Y(G513) );
  NAND2X1 gate135 ( .A(G422), .B(G423), .Y(G516) );
  NAND2X1 gate136 ( .A(G424), .B(G425), .Y(G519) );
  NAND2X1 gate137 ( .A(G426), .B(G429), .Y(G522) );
  NAND2X1 gate138 ( .A(G432), .B(G435), .Y(G525) );
  NAND2X1 gate139 ( .A(G438), .B(G441), .Y(G528) );
  NAND2X1 gate140 ( .A(G444), .B(G447), .Y(G531) );
  NAND2X1 gate141 ( .A(G450), .B(G453), .Y(G534) );
  NAND2X1 gate142 ( .A(G456), .B(G459), .Y(G537) );
  NAND2X1 gate143 ( .A(G462), .B(G465), .Y(G540) );
  NAND2X1 gate144 ( .A(G468), .B(G471), .Y(G543) );
  NAND2X1 gate145 ( .A(G474), .B(G477), .Y(G546) );
  NAND2X1 gate146 ( .A(G480), .B(G483), .Y(G549) );
  NAND2X1 gate147 ( .A(G486), .B(G489), .Y(G552) );
  NAND2X1 gate148 ( .A(G492), .B(G495), .Y(G555) );
  NAND2X1 gate149 ( .A(G498), .B(G501), .Y(G558) );
  NAND2X1 gate150 ( .A(G504), .B(G507), .Y(G561) );
  NAND2X1 gate151 ( .A(G510), .B(G513), .Y(G564) );
  NAND2X1 gate152 ( .A(G516), .B(G519), .Y(G567) );
  NAND2X1 gate153 ( .A(G426), .B(G522), .Y(G570) );
  NAND2X1 gate154 ( .A(G429), .B(G522), .Y(G571) );
  NAND2X1 gate155 ( .A(G432), .B(G525), .Y(G572) );
  NAND2X1 gate156 ( .A(G435), .B(G525), .Y(G573) );
  NAND2X1 gate157 ( .A(G438), .B(G528), .Y(G574) );
  NAND2X1 gate158 ( .A(G441), .B(G528), .Y(G575) );
  NAND2X1 gate159 ( .A(G444), .B(G531), .Y(G576) );
  NAND2X1 gate160 ( .A(G447), .B(G531), .Y(G577) );
  NAND2X1 gate161 ( .A(G450), .B(G534), .Y(G578) );
  NAND2X1 gate162 ( .A(G453), .B(G534), .Y(G579) );
  NAND2X1 gate163 ( .A(G456), .B(G537), .Y(G580) );
  NAND2X1 gate164 ( .A(G459), .B(G537), .Y(G581) );
  NAND2X1 gate165 ( .A(G462), .B(G540), .Y(G582) );
  NAND2X1 gate166 ( .A(G465), .B(G540), .Y(G583) );
  NAND2X1 gate167 ( .A(G468), .B(G543), .Y(G584) );
  NAND2X1 gate168 ( .A(G471), .B(G543), .Y(G585) );
  NAND2X1 gate169 ( .A(G474), .B(G546), .Y(G586) );
  NAND2X1 gate170 ( .A(G477), .B(G546), .Y(G587) );
  NAND2X1 gate171 ( .A(G480), .B(G549), .Y(G588) );
  NAND2X1 gate172 ( .A(G483), .B(G549), .Y(G589) );
  NAND2X1 gate173 ( .A(G486), .B(G552), .Y(G590) );
  NAND2X1 gate174 ( .A(G489), .B(G552), .Y(G591) );
  NAND2X1 gate175 ( .A(G492), .B(G555), .Y(G592) );
  NAND2X1 gate176 ( .A(G495), .B(G555), .Y(G593) );
  NAND2X1 gate177 ( .A(G498), .B(G558), .Y(G594) );
  NAND2X1 gate178 ( .A(G501), .B(G558), .Y(G595) );
  NAND2X1 gate179 ( .A(G504), .B(G561), .Y(G596) );
  NAND2X1 gate180 ( .A(G507), .B(G561), .Y(G597) );
  NAND2X1 gate181 ( .A(G510), .B(G564), .Y(G598) );
  NAND2X1 gate182 ( .A(G513), .B(G564), .Y(G599) );
  NAND2X1 gate183 ( .A(G516), .B(G567), .Y(G600) );
  NAND2X1 gate184 ( .A(G519), .B(G567), .Y(G601) );
  NAND2X1 gate185 ( .A(G570), .B(G571), .Y(G602) );
  NAND2X1 gate186 ( .A(G572), .B(G573), .Y(G607) );
  NAND2X1 gate187 ( .A(G574), .B(G575), .Y(G612) );
  NAND2X1 gate188 ( .A(G576), .B(G577), .Y(G617) );
  NAND2X1 gate189 ( .A(G578), .B(G579), .Y(G622) );
  NAND2X1 gate190 ( .A(G580), .B(G581), .Y(G627) );
  NAND2X1 gate191 ( .A(G582), .B(G583), .Y(G632) );
  NAND2X1 gate192 ( .A(G584), .B(G585), .Y(G637) );
  NAND2X1 gate193 ( .A(G586), .B(G587), .Y(G642) );
  NAND2X1 gate194 ( .A(G588), .B(G589), .Y(G645) );
  NAND2X1 gate195 ( .A(G590), .B(G591), .Y(G648) );
  NAND2X1 gate196 ( .A(G592), .B(G593), .Y(G651) );
  NAND2X1 gate197 ( .A(G594), .B(G595), .Y(G654) );
  NAND2X1 gate198 ( .A(G596), .B(G597), .Y(G657) );
  NAND2X1 gate199 ( .A(G598), .B(G599), .Y(G660) );
  NAND2X1 gate200 ( .A(G600), .B(G601), .Y(G663) );
  NAND2X1 gate201 ( .A(G602), .B(G607), .Y(G666) );
  NAND2X1 gate202 ( .A(G612), .B(G617), .Y(G669) );
  NAND2X1 gate203 ( .A(G602), .B(G612), .Y(G672) );
  NAND2X1 gate204 ( .A(G607), .B(G617), .Y(G675) );
  NAND2X1 gate205 ( .A(G622), .B(G627), .Y(G678) );
  NAND2X1 gate206 ( .A(G632), .B(G637), .Y(G681) );
  NAND2X1 gate207 ( .A(G622), .B(G632), .Y(G684) );
  NAND2X1 gate208 ( .A(G627), .B(G637), .Y(G687) );
  NAND2X1 gate209 ( .A(G602), .B(G666), .Y(G690) );
  NAND2X1 gate210 ( .A(G607), .B(G666), .Y(G691) );
  NAND2X1 gate211 ( .A(G612), .B(G669), .Y(G692) );
  NAND2X1 gate212 ( .A(G617), .B(G669), .Y(G693) );
  NAND2X1 gate213 ( .A(G602), .B(G672), .Y(G694) );
  NAND2X1 gate214 ( .A(G612), .B(G672), .Y(G695) );
  NAND2X1 gate215 ( .A(G607), .B(G675), .Y(G696) );
  NAND2X1 gate216 ( .A(G617), .B(G675), .Y(G697) );
  NAND2X1 gate217 ( .A(G622), .B(G678), .Y(G698) );
  NAND2X1 gate218 ( .A(G627), .B(G678), .Y(G699) );
  NAND2X1 gate219 ( .A(G632), .B(G681), .Y(G700) );
  NAND2X1 gate220 ( .A(G637), .B(G681), .Y(G701) );
  NAND2X1 gate221 ( .A(G622), .B(G684), .Y(G702) );
  NAND2X1 gate222 ( .A(G632), .B(G684), .Y(G703) );
  NAND2X1 gate223 ( .A(G627), .B(G687), .Y(G704) );
  NAND2X1 gate224 ( .A(G637), .B(G687), .Y(G705) );
  NAND2X1 gate225 ( .A(G690), .B(G691), .Y(G706) );
  NAND2X1 gate226 ( .A(G692), .B(G693), .Y(G709) );
  NAND2X1 gate227 ( .A(G694), .B(G695), .Y(G712) );
  NAND2X1 gate228 ( .A(G696), .B(G697), .Y(G715) );
  NAND2X1 gate229 ( .A(G698), .B(G699), .Y(G718) );
  NAND2X1 gate230 ( .A(G700), .B(G701), .Y(G721) );
  NAND2X1 gate231 ( .A(G702), .B(G703), .Y(G724) );
  NAND2X1 gate232 ( .A(G704), .B(G705), .Y(G727) );
  NAND2X1 gate233 ( .A(G242), .B(G718), .Y(G730) );
  NAND2X1 gate234 ( .A(G245), .B(G721), .Y(G733) );
  NAND2X1 gate235 ( .A(G248), .B(G724), .Y(G736) );
  NAND2X1 gate236 ( .A(G251), .B(G727), .Y(G739) );
  NAND2X1 gate237 ( .A(G254), .B(G706), .Y(G742) );
  NAND2X1 gate238 ( .A(G257), .B(G709), .Y(G745) );
  NAND2X1 gate239 ( .A(G260), .B(G712), .Y(G748) );
  NAND2X1 gate240 ( .A(G263), .B(G715), .Y(G751) );
  NAND2X1 gate241 ( .A(G242), .B(G730), .Y(G754) );
  NAND2X1 gate242 ( .A(G718), .B(G730), .Y(G755) );
  NAND2X1 gate243 ( .A(G245), .B(G733), .Y(G756) );
  NAND2X1 gate244 ( .A(G721), .B(G733), .Y(G757) );
  NAND2X1 gate245 ( .A(G248), .B(G736), .Y(G758) );
  NAND2X1 gate246 ( .A(G724), .B(G736), .Y(G759) );
  NAND2X1 gate247 ( .A(G251), .B(G739), .Y(G760) );
  NAND2X1 gate248 ( .A(G727), .B(G739), .Y(G761) );
  NAND2X1 gate249 ( .A(G254), .B(G742), .Y(G762) );
  NAND2X1 gate250 ( .A(G706), .B(G742), .Y(G763) );
  NAND2X1 gate251 ( .A(G257), .B(G745), .Y(G764) );
  NAND2X1 gate252 ( .A(G709), .B(G745), .Y(G765) );
  NAND2X1 gate253 ( .A(G260), .B(G748), .Y(G766) );
  NAND2X1 gate254 ( .A(G712), .B(G748), .Y(G767) );
  NAND2X1 gate255 ( .A(G263), .B(G751), .Y(G768) );
  NAND2X1 gate256 ( .A(G715), .B(G751), .Y(G769) );
  NAND2X1 gate257 ( .A(G754), .B(G755), .Y(G770) );
  NAND2X1 gate258 ( .A(G756), .B(G757), .Y(G773) );
  NAND2X1 gate259 ( .A(G758), .B(G759), .Y(G776) );
  NAND2X1 gate260 ( .A(G760), .B(G761), .Y(G779) );
  NAND2X1 gate261 ( .A(G762), .B(G763), .Y(G782) );
  NAND2X1 gate262 ( .A(G764), .B(G765), .Y(G785) );
  NAND2X1 gate263 ( .A(G766), .B(G767), .Y(G788) );
  NAND2X1 gate264 ( .A(G768), .B(G769), .Y(G791) );
  NAND2X1 gate265 ( .A(G642), .B(G770), .Y(G794) );
  NAND2X1 gate266 ( .A(G645), .B(G773), .Y(G797) );
  NAND2X1 gate267 ( .A(G648), .B(G776), .Y(G800) );
  NAND2X1 gate268 ( .A(G651), .B(G779), .Y(G803) );
  NAND2X1 gate269 ( .A(G654), .B(G782), .Y(G806) );
  NAND2X1 gate270 ( .A(G657), .B(G785), .Y(G809) );
  NAND2X1 gate271 ( .A(G660), .B(G788), .Y(G812) );
  NAND2X1 gate272 ( .A(G663), .B(G791), .Y(G815) );
  NAND2X1 gate273 ( .A(G642), .B(G794), .Y(G818) );
  NAND2X1 gate274 ( .A(G770), .B(G794), .Y(G819) );
  NAND2X1 gate275 ( .A(G645), .B(G797), .Y(G820) );
  NAND2X1 gate276 ( .A(G773), .B(G797), .Y(G821) );
  NAND2X1 gate277 ( .A(G648), .B(G800), .Y(G822) );
  NAND2X1 gate278 ( .A(G776), .B(G800), .Y(G823) );
  NAND2X1 gate279 ( .A(G651), .B(G803), .Y(G824) );
  NAND2X1 gate280 ( .A(G779), .B(G803), .Y(G825) );
  NAND2X1 gate281 ( .A(G654), .B(G806), .Y(G826) );
  NAND2X1 gate282 ( .A(G782), .B(G806), .Y(G827) );
  NAND2X1 gate283 ( .A(G657), .B(G809), .Y(G828) );
  NAND2X1 gate284 ( .A(G785), .B(G809), .Y(G829) );
  NAND2X1 gate285 ( .A(G660), .B(G812), .Y(G830) );
  NAND2X1 gate286 ( .A(G788), .B(G812), .Y(G831) );
  NAND2X1 gate287 ( .A(G663), .B(G815), .Y(G832) );
  NAND2X1 gate288 ( .A(G791), .B(G815), .Y(G833) );
  NAND2X1 gate289 ( .A(G818), .B(G819), .Y(G834) );
  NAND2X1 gate290 ( .A(G820), .B(G821), .Y(G847) );
  NAND2X1 gate291 ( .A(G822), .B(G823), .Y(G860) );
  NAND2X1 gate292 ( .A(G824), .B(G825), .Y(G873) );
  NAND2X1 gate293 ( .A(G828), .B(G829), .Y(G886) );
  NAND2X1 gate294 ( .A(G832), .B(G833), .Y(G899) );
  NAND2X1 gate295 ( .A(G830), .B(G831), .Y(G912) );
  NAND2X1 gate296 ( .A(G826), .B(G827), .Y(G925) );
  INVX1 gate297 ( .A(G834), .Y(G938) );
  INVX1 gate298 ( .A(G847), .Y(G939) );
  INVX1 gate299 ( .A(G860), .Y(G940) );
  INVX1 gate300 ( .A(G834), .Y(G941) );
  INVX1 gate301 ( .A(G847), .Y(G942) );
  INVX1 gate302 ( .A(G873), .Y(G943) );
  INVX1 gate303 ( .A(G834), .Y(G944) );
  INVX1 gate304 ( .A(G860), .Y(G945) );
  INVX1 gate305 ( .A(G873), .Y(G946) );
  INVX1 gate306 ( .A(G847), .Y(G947) );
  INVX1 gate307 ( .A(G860), .Y(G948) );
  INVX1 gate308 ( .A(G873), .Y(G949) );
  INVX1 gate309 ( .A(G886), .Y(G950) );
  INVX1 gate310 ( .A(G899), .Y(G951) );
  INVX1 gate311 ( .A(G886), .Y(G952) );
  INVX1 gate312 ( .A(G912), .Y(G953) );
  INVX1 gate313 ( .A(G925), .Y(G954) );
  INVX1 gate314 ( .A(G899), .Y(G955) );
  INVX1 gate315 ( .A(G925), .Y(G956) );
  INVX1 gate316 ( .A(G912), .Y(G957) );
  INVX1 gate317 ( .A(G925), .Y(G958) );
  INVX1 gate318 ( .A(G886), .Y(G959) );
  INVX1 gate319 ( .A(G912), .Y(G960) );
  INVX1 gate320 ( .A(G925), .Y(G961) );
  INVX1 gate321 ( .A(G886), .Y(G962) );
  INVX1 gate322 ( .A(G899), .Y(G963) );
  INVX1 gate323 ( .A(G925), .Y(G964) );
  INVX1 gate324 ( .A(G912), .Y(G965) );
  INVX1 gate325 ( .A(G899), .Y(G966) );
  INVX1 gate326 ( .A(G886), .Y(G967) );
  INVX1 gate327 ( .A(G912), .Y(G968) );
  INVX1 gate328 ( .A(G899), .Y(G969) );
  INVX1 gate329 ( .A(G847), .Y(G970) );
  INVX1 gate330 ( .A(G873), .Y(G971) );
  INVX1 gate331 ( .A(G847), .Y(G972) );
  INVX1 gate332 ( .A(G860), .Y(G973) );
  INVX1 gate333 ( .A(G834), .Y(G974) );
  INVX1 gate334 ( .A(G873), .Y(G975) );
  INVX1 gate335 ( .A(G834), .Y(G976) );
  INVX1 gate336 ( .A(G860), .Y(G977) );
  AND2X1 gate337_1 ( .A(G938), .B(G939), .Y(G978_1) );
  AND2X1 gate337_2 ( .A(G940), .B(G873), .Y(G978_2) );
  AND2X1 gate337 ( .A(G978_1), .B(G978_2), .Y(G978) );
  AND2X1 gate338_1 ( .A(G941), .B(G942), .Y(G979_1) );
  AND2X1 gate338_2 ( .A(G860), .B(G943), .Y(G979_2) );
  AND2X1 gate338 ( .A(G979_1), .B(G979_2), .Y(G979) );
  AND2X1 gate339_1 ( .A(G944), .B(G847), .Y(G980_1) );
  AND2X1 gate339_2 ( .A(G945), .B(G946), .Y(G980_2) );
  AND2X1 gate339 ( .A(G980_1), .B(G980_2), .Y(G980) );
  AND2X1 gate340_1 ( .A(G834), .B(G947), .Y(G981_1) );
  AND2X1 gate340_2 ( .A(G948), .B(G949), .Y(G981_2) );
  AND2X1 gate340 ( .A(G981_1), .B(G981_2), .Y(G981) );
  AND2X1 gate341_1 ( .A(G958), .B(G959), .Y(G982_1) );
  AND2X1 gate341_2 ( .A(G960), .B(G899), .Y(G982_2) );
  AND2X1 gate341 ( .A(G982_1), .B(G982_2), .Y(G982) );
  AND2X1 gate342_1 ( .A(G961), .B(G962), .Y(G983_1) );
  AND2X1 gate342_2 ( .A(G912), .B(G963), .Y(G983_2) );
  AND2X1 gate342 ( .A(G983_1), .B(G983_2), .Y(G983) );
  AND2X1 gate343_1 ( .A(G964), .B(G886), .Y(G984_1) );
  AND2X1 gate343_2 ( .A(G965), .B(G966), .Y(G984_2) );
  AND2X1 gate343 ( .A(G984_1), .B(G984_2), .Y(G984) );
  AND2X1 gate344_1 ( .A(G925), .B(G967), .Y(G985_1) );
  AND2X1 gate344_2 ( .A(G968), .B(G969), .Y(G985_2) );
  AND2X1 gate344 ( .A(G985_1), .B(G985_2), .Y(G985) );
  OR2X1 gate345_1 ( .A(G978), .B(G979), .Y(G986_1) );
  OR2X1 gate345_2 ( .A(G980), .B(G981), .Y(G986_2) );
  OR2X1 gate345 ( .A(G986_1), .B(G986_2), .Y(G986) );
  OR2X1 gate346_1 ( .A(G982), .B(G983), .Y(G991_1) );
  OR2X1 gate346_2 ( .A(G984), .B(G985), .Y(G991_2) );
  OR2X1 gate346 ( .A(G991_1), .B(G991_2), .Y(G991) );
  AND2X1 gate347_1 ( .A(G925), .B(G950), .Y(G996_1) );
  AND2X1 gate347_2 ( .A(G912), .B(G951), .Y(G996_2) );
  AND2X1 gate347_3 ( .A(G986), .B(G996_1), .Y(G996_3) );
  AND2X1 gate347 ( .A(G996_2), .B(G996_3), .Y(G996) );
  AND2X1 gate348_1 ( .A(G925), .B(G952), .Y(G1001_1) );
  AND2X1 gate348_2 ( .A(G953), .B(G899), .Y(G1001_2) );
  AND2X1 gate348_3 ( .A(G986), .B(G1001_1), .Y(G1001_3) );
  AND2X1 gate348 ( .A(G1001_2), .B(G1001_3), .Y(G1001) );
  AND2X1 gate349_1 ( .A(G954), .B(G886), .Y(G1006_1) );
  AND2X1 gate349_2 ( .A(G912), .B(G955), .Y(G1006_2) );
  AND2X1 gate349_3 ( .A(G986), .B(G1006_1), .Y(G1006_3) );
  AND2X1 gate349 ( .A(G1006_2), .B(G1006_3), .Y(G1006) );
  AND2X1 gate350_1 ( .A(G956), .B(G886), .Y(G1011_1) );
  AND2X1 gate350_2 ( .A(G957), .B(G899), .Y(G1011_2) );
  AND2X1 gate350_3 ( .A(G986), .B(G1011_1), .Y(G1011_3) );
  AND2X1 gate350 ( .A(G1011_2), .B(G1011_3), .Y(G1011) );
  AND2X1 gate351_1 ( .A(G834), .B(G970), .Y(G1016_1) );
  AND2X1 gate351_2 ( .A(G860), .B(G971), .Y(G1016_2) );
  AND2X1 gate351_3 ( .A(G991), .B(G1016_1), .Y(G1016_3) );
  AND2X1 gate351 ( .A(G1016_2), .B(G1016_3), .Y(G1016) );
  AND2X1 gate352_1 ( .A(G834), .B(G972), .Y(G1021_1) );
  AND2X1 gate352_2 ( .A(G973), .B(G873), .Y(G1021_2) );
  AND2X1 gate352_3 ( .A(G991), .B(G1021_1), .Y(G1021_3) );
  AND2X1 gate352 ( .A(G1021_2), .B(G1021_3), .Y(G1021) );
  AND2X1 gate353_1 ( .A(G974), .B(G847), .Y(G1026_1) );
  AND2X1 gate353_2 ( .A(G860), .B(G975), .Y(G1026_2) );
  AND2X1 gate353_3 ( .A(G991), .B(G1026_1), .Y(G1026_3) );
  AND2X1 gate353 ( .A(G1026_2), .B(G1026_3), .Y(G1026) );
  AND2X1 gate354_1 ( .A(G976), .B(G847), .Y(G1031_1) );
  AND2X1 gate354_2 ( .A(G977), .B(G873), .Y(G1031_2) );
  AND2X1 gate354_3 ( .A(G991), .B(G1031_1), .Y(G1031_3) );
  AND2X1 gate354 ( .A(G1031_2), .B(G1031_3), .Y(G1031) );
  AND2X1 gate355 ( .A(G834), .B(G996), .Y(G1036) );
  AND2X1 gate356 ( .A(G847), .B(G996), .Y(G1039) );
  AND2X1 gate357 ( .A(G860), .B(G996), .Y(G1042) );
  AND2X1 gate358 ( .A(G873), .B(G996), .Y(G1045) );
  AND2X1 gate359 ( .A(G834), .B(G1001), .Y(G1048) );
  AND2X1 gate360 ( .A(G847), .B(G1001), .Y(G1051) );
  AND2X1 gate361 ( .A(G860), .B(G1001), .Y(G1054) );
  AND2X1 gate362 ( .A(G873), .B(G1001), .Y(G1057) );
  AND2X1 gate363 ( .A(G834), .B(G1006), .Y(G1060) );
  AND2X1 gate364 ( .A(G847), .B(G1006), .Y(G1063) );
  AND2X1 gate365 ( .A(G860), .B(G1006), .Y(G1066) );
  AND2X1 gate366 ( .A(G873), .B(G1006), .Y(G1069) );
  AND2X1 gate367 ( .A(G834), .B(G1011), .Y(G1072) );
  AND2X1 gate368 ( .A(G847), .B(G1011), .Y(G1075) );
  AND2X1 gate369 ( .A(G860), .B(G1011), .Y(G1078) );
  AND2X1 gate370 ( .A(G873), .B(G1011), .Y(G1081) );
  AND2X1 gate371 ( .A(G925), .B(G1016), .Y(G1084) );
  AND2X1 gate372 ( .A(G886), .B(G1016), .Y(G1087) );
  AND2X1 gate373 ( .A(G912), .B(G1016), .Y(G1090) );
  AND2X1 gate374 ( .A(G899), .B(G1016), .Y(G1093) );
  AND2X1 gate375 ( .A(G925), .B(G1021), .Y(G1096) );
  AND2X1 gate376 ( .A(G886), .B(G1021), .Y(G1099) );
  AND2X1 gate377 ( .A(G912), .B(G1021), .Y(G1102) );
  AND2X1 gate378 ( .A(G899), .B(G1021), .Y(G1105) );
  AND2X1 gate379 ( .A(G925), .B(G1026), .Y(G1108) );
  AND2X1 gate380 ( .A(G886), .B(G1026), .Y(G1111) );
  AND2X1 gate381 ( .A(G912), .B(G1026), .Y(G1114) );
  AND2X1 gate382 ( .A(G899), .B(G1026), .Y(G1117) );
  AND2X1 gate383 ( .A(G925), .B(G1031), .Y(G1120) );
  AND2X1 gate384 ( .A(G886), .B(G1031), .Y(G1123) );
  AND2X1 gate385 ( .A(G912), .B(G1031), .Y(G1126) );
  AND2X1 gate386 ( .A(G899), .B(G1031), .Y(G1129) );
  NAND2X1 gate387 ( .A(G1), .B(G1036), .Y(G1132) );
  NAND2X1 gate388 ( .A(G2), .B(G1039), .Y(G1135) );
  NAND2X1 gate389 ( .A(G3), .B(G1042), .Y(G1138) );
  NAND2X1 gate390 ( .A(G4), .B(G1045), .Y(G1141) );
  NAND2X1 gate391 ( .A(G5), .B(G1048), .Y(G1144) );
  NAND2X1 gate392 ( .A(G6), .B(G1051), .Y(G1147) );
  NAND2X1 gate393 ( .A(G7), .B(G1054), .Y(G1150) );
  NAND2X1 gate394 ( .A(G8), .B(G1057), .Y(G1153) );
  NAND2X1 gate395 ( .A(G9), .B(G1060), .Y(G1156) );
  NAND2X1 gate396 ( .A(G10), .B(G1063), .Y(G1159) );
  NAND2X1 gate397 ( .A(G11), .B(G1066), .Y(G1162) );
  NAND2X1 gate398 ( .A(G12), .B(G1069), .Y(G1165) );
  NAND2X1 gate399 ( .A(G13), .B(G1072), .Y(G1168) );
  NAND2X1 gate400 ( .A(G14), .B(G1075), .Y(G1171) );
  NAND2X1 gate401 ( .A(G15), .B(G1078), .Y(G1174) );
  NAND2X1 gate402 ( .A(G16), .B(G1081), .Y(G1177) );
  NAND2X1 gate403 ( .A(G17), .B(G1084), .Y(G1180) );
  NAND2X1 gate404 ( .A(G18), .B(G1087), .Y(G1183) );
  NAND2X1 gate405 ( .A(G19), .B(G1090), .Y(G1186) );
  NAND2X1 gate406 ( .A(G20), .B(G1093), .Y(G1189) );
  NAND2X1 gate407 ( .A(G21), .B(G1096), .Y(G1192) );
  NAND2X1 gate408 ( .A(G22), .B(G1099), .Y(G1195) );
  NAND2X1 gate409 ( .A(G23), .B(G1102), .Y(G1198) );
  NAND2X1 gate410 ( .A(G24), .B(G1105), .Y(G1201) );
  NAND2X1 gate411 ( .A(G25), .B(G1108), .Y(G1204) );
  NAND2X1 gate412 ( .A(G26), .B(G1111), .Y(G1207) );
  NAND2X1 gate413 ( .A(G27), .B(G1114), .Y(G1210) );
  NAND2X1 gate414 ( .A(G28), .B(G1117), .Y(G1213) );
  NAND2X1 gate415 ( .A(G29), .B(G1120), .Y(G1216) );
  NAND2X1 gate416 ( .A(G30), .B(G1123), .Y(G1219) );
  NAND2X1 gate417 ( .A(G31), .B(G1126), .Y(G1222) );
  NAND2X1 gate418 ( .A(G32), .B(G1129), .Y(G1225) );
  NAND2X1 gate419 ( .A(G1), .B(G1132), .Y(G1228) );
  NAND2X1 gate420 ( .A(G1036), .B(G1132), .Y(G1229) );
  NAND2X1 gate421 ( .A(G2), .B(G1135), .Y(G1230) );
  NAND2X1 gate422 ( .A(G1039), .B(G1135), .Y(G1231) );
  NAND2X1 gate423 ( .A(G3), .B(G1138), .Y(G1232) );
  NAND2X1 gate424 ( .A(G1042), .B(G1138), .Y(G1233) );
  NAND2X1 gate425 ( .A(G4), .B(G1141), .Y(G1234) );
  NAND2X1 gate426 ( .A(G1045), .B(G1141), .Y(G1235) );
  NAND2X1 gate427 ( .A(G5), .B(G1144), .Y(G1236) );
  NAND2X1 gate428 ( .A(G1048), .B(G1144), .Y(G1237) );
  NAND2X1 gate429 ( .A(G6), .B(G1147), .Y(G1238) );
  NAND2X1 gate430 ( .A(G1051), .B(G1147), .Y(G1239) );
  NAND2X1 gate431 ( .A(G7), .B(G1150), .Y(G1240) );
  NAND2X1 gate432 ( .A(G1054), .B(G1150), .Y(G1241) );
  NAND2X1 gate433 ( .A(G8), .B(G1153), .Y(G1242) );
  NAND2X1 gate434 ( .A(G1057), .B(G1153), .Y(G1243) );
  NAND2X1 gate435 ( .A(G9), .B(G1156), .Y(G1244) );
  NAND2X1 gate436 ( .A(G1060), .B(G1156), .Y(G1245) );
  NAND2X1 gate437 ( .A(G10), .B(G1159), .Y(G1246) );
  NAND2X1 gate438 ( .A(G1063), .B(G1159), .Y(G1247) );
  NAND2X1 gate439 ( .A(G11), .B(G1162), .Y(G1248) );
  NAND2X1 gate440 ( .A(G1066), .B(G1162), .Y(G1249) );
  NAND2X1 gate441 ( .A(G12), .B(G1165), .Y(G1250) );
  NAND2X1 gate442 ( .A(G1069), .B(G1165), .Y(G1251) );
  NAND2X1 gate443 ( .A(G13), .B(G1168), .Y(G1252) );
  NAND2X1 gate444 ( .A(G1072), .B(G1168), .Y(G1253) );
  NAND2X1 gate445 ( .A(G14), .B(G1171), .Y(G1254) );
  NAND2X1 gate446 ( .A(G1075), .B(G1171), .Y(G1255) );
  NAND2X1 gate447 ( .A(G15), .B(G1174), .Y(G1256) );
  NAND2X1 gate448 ( .A(G1078), .B(G1174), .Y(G1257) );
  NAND2X1 gate449 ( .A(G16), .B(G1177), .Y(G1258) );
  NAND2X1 gate450 ( .A(G1081), .B(G1177), .Y(G1259) );
  NAND2X1 gate451 ( .A(G17), .B(G1180), .Y(G1260) );
  NAND2X1 gate452 ( .A(G1084), .B(G1180), .Y(G1261) );
  NAND2X1 gate453 ( .A(G18), .B(G1183), .Y(G1262) );
  NAND2X1 gate454 ( .A(G1087), .B(G1183), .Y(G1263) );
  NAND2X1 gate455 ( .A(G19), .B(G1186), .Y(G1264) );
  NAND2X1 gate456 ( .A(G1090), .B(G1186), .Y(G1265) );
  NAND2X1 gate457 ( .A(G20), .B(G1189), .Y(G1266) );
  NAND2X1 gate458 ( .A(G1093), .B(G1189), .Y(G1267) );
  NAND2X1 gate459 ( .A(G21), .B(G1192), .Y(G1268) );
  NAND2X1 gate460 ( .A(G1096), .B(G1192), .Y(G1269) );
  NAND2X1 gate461 ( .A(G22), .B(G1195), .Y(G1270) );
  NAND2X1 gate462 ( .A(G1099), .B(G1195), .Y(G1271) );
  NAND2X1 gate463 ( .A(G23), .B(G1198), .Y(G1272) );
  NAND2X1 gate464 ( .A(G1102), .B(G1198), .Y(G1273) );
  NAND2X1 gate465 ( .A(G24), .B(G1201), .Y(G1274) );
  NAND2X1 gate466 ( .A(G1105), .B(G1201), .Y(G1275) );
  NAND2X1 gate467 ( .A(G25), .B(G1204), .Y(G1276) );
  NAND2X1 gate468 ( .A(G1108), .B(G1204), .Y(G1277) );
  NAND2X1 gate469 ( .A(G26), .B(G1207), .Y(G1278) );
  NAND2X1 gate470 ( .A(G1111), .B(G1207), .Y(G1279) );
  NAND2X1 gate471 ( .A(G27), .B(G1210), .Y(G1280) );
  NAND2X1 gate472 ( .A(G1114), .B(G1210), .Y(G1281) );
  NAND2X1 gate473 ( .A(G28), .B(G1213), .Y(G1282) );
  NAND2X1 gate474 ( .A(G1117), .B(G1213), .Y(G1283) );
  NAND2X1 gate475 ( .A(G29), .B(G1216), .Y(G1284) );
  NAND2X1 gate476 ( .A(G1120), .B(G1216), .Y(G1285) );
  NAND2X1 gate477 ( .A(G30), .B(G1219), .Y(G1286) );
  NAND2X1 gate478 ( .A(G1123), .B(G1219), .Y(G1287) );
  NAND2X1 gate479 ( .A(G31), .B(G1222), .Y(G1288) );
  NAND2X1 gate480 ( .A(G1126), .B(G1222), .Y(G1289) );
  NAND2X1 gate481 ( .A(G32), .B(G1225), .Y(G1290) );
  NAND2X1 gate482 ( .A(G1129), .B(G1225), .Y(G1291) );
  NAND2X1 gate483 ( .A(G1228), .B(G1229), .Y(G1292) );
  NAND2X1 gate484 ( .A(G1230), .B(G1231), .Y(G1293) );
  NAND2X1 gate485 ( .A(G1232), .B(G1233), .Y(G1294) );
  NAND2X1 gate486 ( .A(G1234), .B(G1235), .Y(G1295) );
  NAND2X1 gate487 ( .A(G1236), .B(G1237), .Y(G1296) );
  NAND2X1 gate488 ( .A(G1238), .B(G1239), .Y(G1297) );
  NAND2X1 gate489 ( .A(G1240), .B(G1241), .Y(G1298) );
  NAND2X1 gate490 ( .A(G1242), .B(G1243), .Y(G1299) );
  NAND2X1 gate491 ( .A(G1244), .B(G1245), .Y(G1300) );
  NAND2X1 gate492 ( .A(G1246), .B(G1247), .Y(G1301) );
  NAND2X1 gate493 ( .A(G1248), .B(G1249), .Y(G1302) );
  NAND2X1 gate494 ( .A(G1250), .B(G1251), .Y(G1303) );
  NAND2X1 gate495 ( .A(G1252), .B(G1253), .Y(G1304) );
  NAND2X1 gate496 ( .A(G1254), .B(G1255), .Y(G1305) );
  NAND2X1 gate497 ( .A(G1256), .B(G1257), .Y(G1306) );
  NAND2X1 gate498 ( .A(G1258), .B(G1259), .Y(G1307) );
  NAND2X1 gate499 ( .A(G1260), .B(G1261), .Y(G1308) );
  NAND2X1 gate500 ( .A(G1262), .B(G1263), .Y(G1309) );
  NAND2X1 gate501 ( .A(G1264), .B(G1265), .Y(G1310) );
  NAND2X1 gate502 ( .A(G1266), .B(G1267), .Y(G1311) );
  NAND2X1 gate503 ( .A(G1268), .B(G1269), .Y(G1312) );
  NAND2X1 gate504 ( .A(G1270), .B(G1271), .Y(G1313) );
  NAND2X1 gate505 ( .A(G1272), .B(G1273), .Y(G1314) );
  NAND2X1 gate506 ( .A(G1274), .B(G1275), .Y(G1315) );
  NAND2X1 gate507 ( .A(G1276), .B(G1277), .Y(G1316) );
  NAND2X1 gate508 ( .A(G1278), .B(G1279), .Y(G1317) );
  NAND2X1 gate509 ( .A(G1280), .B(G1281), .Y(G1318) );
  NAND2X1 gate510 ( .A(G1282), .B(G1283), .Y(G1319) );
  NAND2X1 gate511 ( .A(G1284), .B(G1285), .Y(G1320) );
  NAND2X1 gate512 ( .A(G1286), .B(G1287), .Y(G1321) );
  NAND2X1 gate513 ( .A(G1288), .B(G1289), .Y(G1322) );
  NAND2X1 gate514 ( .A(G1290), .B(G1291), .Y(G1323) );
  INVX1 gate515 ( .A(G1292), .Y(G1324) );
  INVX1 gate516 ( .A(G1293), .Y(G1325) );
  INVX1 gate517 ( .A(G1294), .Y(G1326) );
  INVX1 gate518 ( .A(G1295), .Y(G1327) );
  INVX1 gate519 ( .A(G1296), .Y(G1328) );
  INVX1 gate520 ( .A(G1297), .Y(G1329) );
  INVX1 gate521 ( .A(G1298), .Y(G1330) );
  INVX1 gate522 ( .A(G1299), .Y(G1331) );
  INVX1 gate523 ( .A(G1300), .Y(G1332) );
  INVX1 gate524 ( .A(G1301), .Y(G1333) );
  INVX1 gate525 ( .A(G1302), .Y(G1334) );
  INVX1 gate526 ( .A(G1303), .Y(G1335) );
  INVX1 gate527 ( .A(G1304), .Y(G1336) );
  INVX1 gate528 ( .A(G1305), .Y(G1337) );
  INVX1 gate529 ( .A(G1306), .Y(G1338) );
  INVX1 gate530 ( .A(G1307), .Y(G1339) );
  INVX1 gate531 ( .A(G1308), .Y(G1340) );
  INVX1 gate532 ( .A(G1309), .Y(G1341) );
  INVX1 gate533 ( .A(G1310), .Y(G1342) );
  INVX1 gate534 ( .A(G1311), .Y(G1343) );
  INVX1 gate535 ( .A(G1312), .Y(G1344) );
  INVX1 gate536 ( .A(G1313), .Y(G1345) );
  INVX1 gate537 ( .A(G1314), .Y(G1346) );
  INVX1 gate538 ( .A(G1315), .Y(G1347) );
  INVX1 gate539 ( .A(G1316), .Y(G1348) );
  INVX1 gate540 ( .A(G1317), .Y(G1349) );
  INVX1 gate541 ( .A(G1318), .Y(G1350) );
  INVX1 gate542 ( .A(G1319), .Y(G1351) );
  INVX1 gate543 ( .A(G1320), .Y(G1352) );
  INVX1 gate544 ( .A(G1321), .Y(G1353) );
  INVX1 gate545 ( .A(G1322), .Y(G1354) );
  INVX1 gate546 ( .A(G1323), .Y(G1355) );
endmodule


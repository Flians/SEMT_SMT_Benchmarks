
module c6288_synth ( N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, 
        N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, 
        N392, N409, N426, N443, N460, N477, N494, N511, N528, N545, N1581, 
        N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, 
        N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, 
        N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288
 );
  input N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205,
         N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392,
         N409, N426, N443, N460, N477, N494, N511, N528;
  output N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241,
         N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180,
         N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280,
         N6287, N6288;
  wire   N546, N549, N552, N555, N558, N561, N564, N567, N570, N573, N576,
         N579, N582, N585, N588, N591, N594, N597, N600, N603, N606, N609,
         N612, N615, N618, N621, N624, N627, N630, N633, N636, N639, N642,
         N645, N648, N651, N654, N657, N660, N663, N666, N669, N672, N675,
         N678, N681, N684, N687, N690, N693, N696, N699, N702, N705, N708,
         N711, N714, N717, N720, N723, N726, N729, N732, N735, N738, N741,
         N744, N747, N750, N753, N756, N759, N762, N765, N768, N771, N774,
         N777, N780, N783, N786, N789, N792, N795, N798, N801, N804, N807,
         N810, N813, N816, N819, N822, N825, N828, N831, N834, N837, N840,
         N843, N846, N849, N852, N855, N858, N861, N864, N867, N870, N873,
         N876, N879, N882, N885, N888, N891, N894, N897, N900, N903, N906,
         N909, N912, N915, N918, N921, N924, N927, N930, N933, N936, N939,
         N942, N945, N948, N951, N954, N957, N960, N963, N966, N969, N972,
         N975, N978, N981, N984, N987, N990, N993, N996, N999, N1002, N1005,
         N1008, N1011, N1014, N1017, N1020, N1023, N1026, N1029, N1032, N1035,
         N1038, N1041, N1044, N1047, N1050, N1053, N1056, N1059, N1062, N1065,
         N1068, N1071, N1074, N1077, N1080, N1083, N1086, N1089, N1092, N1095,
         N1098, N1101, N1104, N1107, N1110, N1113, N1116, N1119, N1122, N1125,
         N1128, N1131, N1134, N1137, N1140, N1143, N1146, N1149, N1152, N1155,
         N1158, N1161, N1164, N1167, N1170, N1173, N1176, N1179, N1182, N1185,
         N1188, N1191, N1194, N1197, N1200, N1203, N1206, N1209, N1212, N1215,
         N1218, N1221, N1224, N1227, N1230, N1233, N1236, N1239, N1242, N1245,
         N1248, N1251, N1254, N1257, N1260, N1263, N1266, N1269, N1272, N1275,
         N1278, N1281, N1284, N1287, N1290, N1293, N1296, N1299, N1302, N1305,
         N1308, N1311, N1315, N1319, N1323, N1327, N1331, N1335, N1339, N1343,
         N1347, N1351, N1355, N1359, N1363, N1367, N1371, N1372, N1373, N1374,
         N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384,
         N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394,
         N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1404, N1407, N1410,
         N1413, N1416, N1419, N1422, N1425, N1428, N1431, N1434, N1437, N1440,
         N1443, N1446, N1450, N1454, N1458, N1462, N1466, N1470, N1474, N1478,
         N1482, N1486, N1490, N1494, N1498, N1502, N1506, N1507, N1508, N1511,
         N1512, N1513, N1516, N1517, N1518, N1521, N1522, N1523, N1526, N1527,
         N1528, N1531, N1532, N1533, N1536, N1537, N1538, N1541, N1542, N1543,
         N1546, N1547, N1548, N1551, N1552, N1553, N1556, N1557, N1558, N1561,
         N1562, N1563, N1566, N1567, N1568, N1571, N1572, N1573, N1576, N1577,
         N1578, N1582, N1585, N1588, N1591, N1594, N1597, N1600, N1603, N1606,
         N1609, N1612, N1615, N1618, N1621, N1624, N1628, N1632, N1636, N1640,
         N1644, N1648, N1652, N1656, N1660, N1664, N1668, N1672, N1676, N1680,
         N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692, N1693,
         N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702, N1703,
         N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712, N1713,
         N1714, N1717, N1720, N1723, N1726, N1729, N1732, N1735, N1738, N1741,
         N1744, N1747, N1750, N1753, N1756, N1759, N1763, N1767, N1771, N1775,
         N1779, N1783, N1787, N1791, N1795, N1799, N1803, N1807, N1811, N1815,
         N1819, N1820, N1821, N1824, N1825, N1826, N1829, N1830, N1831, N1834,
         N1835, N1836, N1839, N1840, N1841, N1844, N1845, N1846, N1849, N1850,
         N1851, N1854, N1855, N1856, N1859, N1860, N1861, N1864, N1865, N1866,
         N1869, N1870, N1871, N1874, N1875, N1876, N1879, N1880, N1881, N1884,
         N1885, N1886, N1889, N1890, N1891, N1894, N1897, N1902, N1905, N1908,
         N1911, N1914, N1917, N1920, N1923, N1926, N1929, N1932, N1935, N1938,
         N1941, N1945, N1946, N1947, N1951, N1955, N1959, N1963, N1967, N1971,
         N1975, N1979, N1983, N1987, N1991, N1995, N1999, N2000, N2001, N2004,
         N2005, N2006, N2007, N2008, N2009, N2010, N2011, N2012, N2013, N2014,
         N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024,
         N2025, N2026, N2027, N2028, N2029, N2030, N2033, N2037, N2040, N2043,
         N2046, N2049, N2052, N2055, N2058, N2061, N2064, N2067, N2070, N2073,
         N2076, N2080, N2081, N2082, N2085, N2089, N2093, N2097, N2101, N2105,
         N2109, N2113, N2117, N2121, N2125, N2129, N2133, N2137, N2138, N2139,
         N2142, N2145, N2149, N2150, N2151, N2154, N2155, N2156, N2159, N2160,
         N2161, N2164, N2165, N2166, N2169, N2170, N2171, N2174, N2175, N2176,
         N2179, N2180, N2181, N2184, N2185, N2186, N2189, N2190, N2191, N2194,
         N2195, N2196, N2199, N2200, N2201, N2204, N2205, N2206, N2209, N2210,
         N2211, N2214, N2217, N2221, N2222, N2224, N2227, N2230, N2233, N2236,
         N2239, N2242, N2245, N2248, N2251, N2254, N2257, N2260, N2264, N2265,
         N2266, N2269, N2273, N2277, N2281, N2285, N2289, N2293, N2297, N2301,
         N2305, N2309, N2313, N2317, N2318, N2319, N2322, N2326, N2327, N2328,
         N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338,
         N2339, N2340, N2341, N2342, N2343, N2344, N2345, N2346, N2347, N2348,
         N2349, N2350, N2353, N2357, N2358, N2359, N2362, N2365, N2368, N2371,
         N2374, N2377, N2380, N2383, N2386, N2389, N2392, N2395, N2398, N2402,
         N2403, N2404, N2407, N2410, N2414, N2418, N2422, N2426, N2430, N2434,
         N2438, N2442, N2446, N2450, N2454, N2458, N2462, N2463, N2464, N2467,
         N2470, N2474, N2475, N2476, N2477, N2478, N2481, N2482, N2483, N2486,
         N2487, N2488, N2491, N2492, N2493, N2496, N2497, N2498, N2501, N2502,
         N2503, N2506, N2507, N2508, N2511, N2512, N2513, N2516, N2517, N2518,
         N2521, N2522, N2523, N2526, N2527, N2528, N2531, N2532, N2533, N2536,
         N2539, N2543, N2544, N2545, N2549, N2552, N2555, N2558, N2561, N2564,
         N2567, N2570, N2573, N2576, N2579, N2582, N2586, N2587, N2588, N2591,
         N2595, N2599, N2603, N2607, N2611, N2615, N2619, N2623, N2627, N2631,
         N2635, N2639, N2640, N2641, N2644, N2648, N2649, N2650, N2653, N2654,
         N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662, N2663, N2664,
         N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674,
         N2675, N2678, N2682, N2683, N2684, N2687, N2690, N2694, N2697, N2700,
         N2703, N2706, N2709, N2712, N2715, N2718, N2721, N2724, N2727, N2731,
         N2732, N2733, N2736, N2739, N2743, N2744, N2745, N2749, N2753, N2757,
         N2761, N2765, N2769, N2773, N2777, N2781, N2785, N2789, N2790, N2791,
         N2794, N2797, N2801, N2802, N2803, N2806, N2807, N2808, N2811, N2812,
         N2813, N2816, N2817, N2818, N2821, N2822, N2823, N2826, N2827, N2828,
         N2831, N2832, N2833, N2836, N2837, N2838, N2841, N2842, N2843, N2846,
         N2847, N2848, N2851, N2852, N2853, N2856, N2857, N2858, N2861, N2864,
         N2868, N2869, N2870, N2873, N2878, N2881, N2884, N2887, N2890, N2893,
         N2896, N2899, N2902, N2905, N2908, N2912, N2913, N2914, N2917, N2921,
         N2922, N2923, N2926, N2930, N2934, N2938, N2942, N2946, N2950, N2954,
         N2958, N2962, N2966, N2967, N2968, N2971, N2975, N2976, N2977, N2980,
         N2983, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995,
         N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005,
         N3006, N3007, N3010, N3014, N3015, N3016, N3019, N3022, N3026, N3027,
         N3028, N3031, N3034, N3037, N3040, N3043, N3046, N3049, N3052, N3055,
         N3058, N3062, N3063, N3064, N3067, N3070, N3074, N3075, N3076, N3079,
         N3083, N3087, N3091, N3095, N3099, N3103, N3107, N3111, N3115, N3119,
         N3120, N3121, N3124, N3127, N3131, N3132, N3133, N3136, N3140, N3141,
         N3142, N3145, N3146, N3147, N3150, N3151, N3152, N3155, N3156, N3157,
         N3160, N3161, N3162, N3165, N3166, N3167, N3170, N3171, N3172, N3175,
         N3176, N3177, N3180, N3181, N3182, N3185, N3186, N3187, N3190, N3193,
         N3197, N3198, N3199, N3202, N3206, N3207, N3208, N3212, N3215, N3218,
         N3221, N3224, N3227, N3230, N3233, N3236, N3239, N3243, N3244, N3245,
         N3248, N3252, N3253, N3254, N3257, N3260, N3264, N3268, N3272, N3276,
         N3280, N3284, N3288, N3292, N3296, N3300, N3301, N3302, N3305, N3309,
         N3310, N3311, N3314, N3317, N3321, N3322, N3323, N3324, N3325, N3326,
         N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336,
         N3337, N3338, N3339, N3340, N3341, N3344, N3348, N3349, N3350, N3353,
         N3356, N3360, N3361, N3362, N3365, N3368, N3371, N3374, N3377, N3380,
         N3383, N3386, N3389, N3392, N3396, N3397, N3398, N3401, N3404, N3408,
         N3409, N3410, N3413, N3417, N3421, N3425, N3429, N3433, N3437, N3441,
         N3445, N3449, N3453, N3454, N3455, N3458, N3461, N3465, N3466, N3467,
         N3470, N3474, N3475, N3476, N3479, N3480, N3481, N3484, N3485, N3486,
         N3489, N3490, N3491, N3494, N3495, N3496, N3499, N3500, N3501, N3504,
         N3505, N3506, N3509, N3510, N3511, N3514, N3515, N3516, N3519, N3520,
         N3521, N3524, N3527, N3531, N3532, N3533, N3536, N3540, N3541, N3542,
         N3545, N3548, N3553, N3556, N3559, N3562, N3565, N3568, N3571, N3574,
         N3577, N3581, N3582, N3583, N3586, N3590, N3591, N3592, N3595, N3598,
         N3602, N3603, N3604, N3608, N3612, N3616, N3620, N3624, N3628, N3632,
         N3636, N3637, N3638, N3641, N3645, N3646, N3647, N3650, N3653, N3657,
         N3658, N3659, N3662, N3663, N3664, N3665, N3666, N3667, N3668, N3669,
         N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3681,
         N3685, N3686, N3687, N3690, N3693, N3697, N3698, N3699, N3702, N3706,
         N3709, N3712, N3715, N3718, N3721, N3724, N3727, N3730, N3734, N3735,
         N3736, N3739, N3742, N3746, N3747, N3748, N3751, N3755, N3756, N3757,
         N3760, N3764, N3768, N3772, N3776, N3780, N3784, N3788, N3792, N3793,
         N3794, N3797, N3800, N3804, N3805, N3806, N3809, N3813, N3814, N3815,
         N3818, N3821, N3825, N3826, N3827, N3830, N3831, N3832, N3835, N3836,
         N3837, N3840, N3841, N3842, N3845, N3846, N3847, N3850, N3851, N3852,
         N3855, N3856, N3857, N3860, N3861, N3862, N3865, N3868, N3872, N3873,
         N3874, N3877, N3881, N3882, N3883, N3886, N3889, N3893, N3894, N3896,
         N3899, N3902, N3905, N3908, N3911, N3914, N3917, N3921, N3922, N3923,
         N3926, N3930, N3931, N3932, N3935, N3938, N3942, N3943, N3944, N3947,
         N3951, N3955, N3959, N3963, N3967, N3971, N3975, N3976, N3977, N3980,
         N3984, N3985, N3986, N3989, N3992, N3996, N3997, N3998, N4001, N4005,
         N4006, N4007, N4008, N4009, N4010, N4011, N4012, N4013, N4014, N4015,
         N4016, N4017, N4018, N4019, N4022, N4026, N4027, N4028, N4031, N4034,
         N4038, N4039, N4040, N4043, N4047, N4048, N4049, N4052, N4055, N4058,
         N4061, N4064, N4067, N4070, N4073, N4077, N4078, N4079, N4082, N4085,
         N4089, N4090, N4091, N4094, N4098, N4099, N4100, N4103, N4106, N4110,
         N4114, N4118, N4122, N4126, N4130, N4134, N4138, N4139, N4140, N4143,
         N4146, N4150, N4151, N4152, N4155, N4159, N4160, N4161, N4164, N4167,
         N4171, N4172, N4173, N4174, N4175, N4178, N4179, N4180, N4183, N4184,
         N4185, N4188, N4189, N4190, N4193, N4194, N4195, N4198, N4199, N4200,
         N4203, N4204, N4205, N4208, N4211, N4215, N4216, N4217, N4220, N4224,
         N4225, N4226, N4229, N4232, N4236, N4237, N4238, N4242, N4245, N4248,
         N4251, N4254, N4257, N4260, N4264, N4265, N4266, N4269, N4273, N4274,
         N4275, N4278, N4281, N4285, N4286, N4287, N4290, N4294, N4298, N4302,
         N4306, N4310, N4314, N4318, N4319, N4320, N4323, N4327, N4328, N4329,
         N4332, N4335, N4339, N4340, N4341, N4344, N4348, N4349, N4350, N4353,
         N4354, N4355, N4356, N4357, N4358, N4359, N4360, N4361, N4362, N4363,
         N4364, N4365, N4368, N4372, N4373, N4374, N4377, N4380, N4384, N4385,
         N4386, N4389, N4393, N4394, N4395, N4398, N4401, N4405, N4408, N4411,
         N4414, N4417, N4420, N4423, N4427, N4428, N4429, N4432, N4435, N4439,
         N4440, N4441, N4444, N4448, N4449, N4450, N4453, N4456, N4460, N4461,
         N4462, N4466, N4470, N4474, N4478, N4482, N4486, N4487, N4488, N4491,
         N4494, N4498, N4499, N4500, N4503, N4507, N4508, N4509, N4512, N4515,
         N4519, N4520, N4521, N4524, N4525, N4526, N4529, N4530, N4531, N4534,
         N4535, N4536, N4539, N4540, N4541, N4544, N4545, N4546, N4549, N4550,
         N4551, N4554, N4557, N4561, N4562, N4563, N4566, N4570, N4571, N4572,
         N4575, N4578, N4582, N4583, N4584, N4587, N4592, N4595, N4598, N4601,
         N4604, N4607, N4611, N4612, N4613, N4616, N4620, N4621, N4622, N4625,
         N4628, N4632, N4633, N4634, N4637, N4641, N4642, N4643, N4646, N4650,
         N4654, N4658, N4662, N4666, N4667, N4668, N4671, N4675, N4676, N4677,
         N4680, N4683, N4687, N4688, N4689, N4692, N4696, N4697, N4698, N4701,
         N4704, N4708, N4709, N4710, N4711, N4712, N4713, N4714, N4715, N4716,
         N4717, N4718, N4721, N4725, N4726, N4727, N4730, N4733, N4737, N4738,
         N4739, N4742, N4746, N4747, N4748, N4751, N4754, N4758, N4759, N4760,
         N4763, N4766, N4769, N4772, N4775, N4779, N4780, N4781, N4784, N4787,
         N4791, N4792, N4793, N4796, N4800, N4801, N4802, N4805, N4808, N4812,
         N4813, N4814, N4817, N4821, N4825, N4829, N4833, N4837, N4838, N4839,
         N4842, N4845, N4849, N4850, N4851, N4854, N4858, N4859, N4860, N4863,
         N4866, N4870, N4871, N4872, N4875, N4879, N4880, N4881, N4884, N4885,
         N4886, N4889, N4890, N4891, N4894, N4895, N4896, N4899, N4900, N4901,
         N4904, N4907, N4911, N4912, N4913, N4916, N4920, N4921, N4922, N4925,
         N4928, N4932, N4933, N4934, N4937, N4941, N4942, N4943, N4947, N4950,
         N4953, N4956, N4959, N4963, N4964, N4965, N4968, N4972, N4973, N4974,
         N4977, N4980, N4984, N4985, N4986, N4989, N4993, N4994, N4995, N4998,
         N5001, N5005, N5009, N5013, N5017, N5021, N5022, N5023, N5026, N5030,
         N5031, N5032, N5035, N5038, N5042, N5043, N5044, N5047, N5051, N5052,
         N5053, N5056, N5059, N5063, N5064, N5065, N5066, N5067, N5068, N5069,
         N5070, N5071, N5072, N5073, N5076, N5080, N5081, N5082, N5085, N5088,
         N5092, N5093, N5094, N5097, N5101, N5102, N5103, N5106, N5109, N5113,
         N5114, N5115, N5118, N5121, N5124, N5127, N5130, N5134, N5135, N5136,
         N5139, N5142, N5146, N5147, N5148, N5151, N5155, N5156, N5157, N5160,
         N5163, N5167, N5168, N5169, N5172, N5176, N5180, N5184, N5188, N5192,
         N5193, N5194, N5197, N5200, N5204, N5205, N5206, N5209, N5213, N5214,
         N5215, N5218, N5221, N5225, N5226, N5227, N5230, N5234, N5235, N5236,
         N5239, N5240, N5241, N5244, N5245, N5246, N5249, N5250, N5251, N5254,
         N5255, N5256, N5259, N5262, N5266, N5267, N5268, N5271, N5275, N5276,
         N5277, N5280, N5283, N5287, N5288, N5289, N5292, N5296, N5297, N5298,
         N5301, N5304, N5309, N5312, N5315, N5318, N5322, N5323, N5324, N5327,
         N5331, N5332, N5333, N5336, N5339, N5343, N5344, N5345, N5348, N5352,
         N5353, N5354, N5357, N5360, N5364, N5365, N5366, N5370, N5374, N5378,
         N5379, N5380, N5383, N5387, N5388, N5389, N5392, N5395, N5399, N5400,
         N5401, N5404, N5408, N5409, N5410, N5413, N5416, N5420, N5421, N5422,
         N5425, N5426, N5427, N5428, N5429, N5430, N5431, N5434, N5438, N5439,
         N5440, N5443, N5446, N5450, N5451, N5452, N5455, N5459, N5460, N5461,
         N5464, N5467, N5471, N5472, N5473, N5476, N5480, N5483, N5486, N5489,
         N5493, N5494, N5495, N5498, N5501, N5505, N5506, N5507, N5510, N5514,
         N5515, N5516, N5519, N5522, N5526, N5527, N5528, N5531, N5535, N5536,
         N5537, N5540, N5544, N5548, N5552, N5553, N5554, N5557, N5560, N5564,
         N5565, N5566, N5569, N5573, N5574, N5575, N5578, N5581, N5585, N5586,
         N5587, N5590, N5594, N5595, N5596, N5599, N5602, N5606, N5607, N5608,
         N5611, N5612, N5613, N5616, N5617, N5618, N5621, N5624, N5628, N5629,
         N5630, N5633, N5637, N5638, N5639, N5642, N5645, N5649, N5650, N5651,
         N5654, N5658, N5659, N5660, N5663, N5666, N5670, N5671, N5673, N5676,
         N5679, N5683, N5684, N5685, N5688, N5692, N5693, N5694, N5697, N5700,
         N5704, N5705, N5706, N5709, N5713, N5714, N5715, N5718, N5721, N5725,
         N5726, N5727, N5730, N5734, N5738, N5739, N5740, N5743, N5747, N5748,
         N5749, N5752, N5755, N5759, N5760, N5761, N5764, N5768, N5769, N5770,
         N5773, N5776, N5780, N5781, N5782, N5785, N5786, N5787, N5788, N5789,
         N5792, N5796, N5797, N5798, N5801, N5804, N5808, N5809, N5810, N5813,
         N5817, N5818, N5819, N5822, N5825, N5829, N5830, N5831, N5834, N5837,
         N5840, N5844, N5845, N5846, N5849, N5852, N5856, N5857, N5858, N5861,
         N5865, N5866, N5867, N5870, N5873, N5877, N5878, N5879, N5882, N5886,
         N5890, N5891, N5892, N5895, N5898, N5902, N5903, N5904, N5907, N5911,
         N5912, N5913, N5916, N5919, N5923, N5924, N5925, N5928, N5929, N5930,
         N5933, N5934, N5935, N5938, N5941, N5945, N5946, N5947, N5950, N5954,
         N5955, N5956, N5959, N5962, N5966, N5967, N5968, N5972, N5975, N5979,
         N5980, N5981, N5984, N5988, N5989, N5990, N5993, N5996, N6000, N6001,
         N6002, N6005, N6009, N6010, N6011, N6014, N6018, N6019, N6020, N6023,
         N6026, N6030, N6031, N6032, N6035, N6036, N6037, N6040, N6044, N6045,
         N6046, N6049, N6052, N6056, N6057, N6058, N6061, N6064, N6068, N6069,
         N6070, N6073, N6076, N6080, N6081, N6082, N6085, N6089, N6090, N6091,
         N6094, N6097, N6101, N6102, N6103, N6106, N6107, N6108, N6111, N6114,
         N6118, N6119, N6120, N6124, N6128, N6129, N6130, N6133, N6134, N6135,
         N6138, N6141, N6145, N6146, N6147, N6151, N6155, N6156, N6157, N6161,
         N6165, N6166, N6167, N6171, N6175, N6176, N6177, N6181, N6185, N6186,
         N6187, N6191, N6195, N6196, N6197, N6201, N6205, N6206, N6207, N6211,
         N6215, N6216, N6217, N6221, N6225, N6226, N6227, N6231, N6235, N6236,
         N6237, N6241, N6245, N6246, N6247, N6251, N6255, N6256, N6257, N6261,
         N6265, N6266, N6267, N6271, N6275, N6276, N6277, N6281, N6285, N6286;

  AND2X1 gate1 ( .A(N1), .B(N273), .Y(N545) );
  AND2X1 gate2 ( .A(N1), .B(N290), .Y(N546) );
  AND2X1 gate3 ( .A(N1), .B(N307), .Y(N549) );
  AND2X1 gate4 ( .A(N1), .B(N324), .Y(N552) );
  AND2X1 gate5 ( .A(N1), .B(N341), .Y(N555) );
  AND2X1 gate6 ( .A(N1), .B(N358), .Y(N558) );
  AND2X1 gate7 ( .A(N1), .B(N375), .Y(N561) );
  AND2X1 gate8 ( .A(N1), .B(N392), .Y(N564) );
  AND2X1 gate9 ( .A(N1), .B(N409), .Y(N567) );
  AND2X1 gate10 ( .A(N1), .B(N426), .Y(N570) );
  AND2X1 gate11 ( .A(N1), .B(N443), .Y(N573) );
  AND2X1 gate12 ( .A(N1), .B(N460), .Y(N576) );
  AND2X1 gate13 ( .A(N1), .B(N477), .Y(N579) );
  AND2X1 gate14 ( .A(N1), .B(N494), .Y(N582) );
  AND2X1 gate15 ( .A(N1), .B(N511), .Y(N585) );
  AND2X1 gate16 ( .A(N1), .B(N528), .Y(N588) );
  AND2X1 gate17 ( .A(N18), .B(N273), .Y(N591) );
  AND2X1 gate18 ( .A(N18), .B(N290), .Y(N594) );
  AND2X1 gate19 ( .A(N18), .B(N307), .Y(N597) );
  AND2X1 gate20 ( .A(N18), .B(N324), .Y(N600) );
  AND2X1 gate21 ( .A(N18), .B(N341), .Y(N603) );
  AND2X1 gate22 ( .A(N18), .B(N358), .Y(N606) );
  AND2X1 gate23 ( .A(N18), .B(N375), .Y(N609) );
  AND2X1 gate24 ( .A(N18), .B(N392), .Y(N612) );
  AND2X1 gate25 ( .A(N18), .B(N409), .Y(N615) );
  AND2X1 gate26 ( .A(N18), .B(N426), .Y(N618) );
  AND2X1 gate27 ( .A(N18), .B(N443), .Y(N621) );
  AND2X1 gate28 ( .A(N18), .B(N460), .Y(N624) );
  AND2X1 gate29 ( .A(N18), .B(N477), .Y(N627) );
  AND2X1 gate30 ( .A(N18), .B(N494), .Y(N630) );
  AND2X1 gate31 ( .A(N18), .B(N511), .Y(N633) );
  AND2X1 gate32 ( .A(N18), .B(N528), .Y(N636) );
  AND2X1 gate33 ( .A(N35), .B(N273), .Y(N639) );
  AND2X1 gate34 ( .A(N35), .B(N290), .Y(N642) );
  AND2X1 gate35 ( .A(N35), .B(N307), .Y(N645) );
  AND2X1 gate36 ( .A(N35), .B(N324), .Y(N648) );
  AND2X1 gate37 ( .A(N35), .B(N341), .Y(N651) );
  AND2X1 gate38 ( .A(N35), .B(N358), .Y(N654) );
  AND2X1 gate39 ( .A(N35), .B(N375), .Y(N657) );
  AND2X1 gate40 ( .A(N35), .B(N392), .Y(N660) );
  AND2X1 gate41 ( .A(N35), .B(N409), .Y(N663) );
  AND2X1 gate42 ( .A(N35), .B(N426), .Y(N666) );
  AND2X1 gate43 ( .A(N35), .B(N443), .Y(N669) );
  AND2X1 gate44 ( .A(N35), .B(N460), .Y(N672) );
  AND2X1 gate45 ( .A(N35), .B(N477), .Y(N675) );
  AND2X1 gate46 ( .A(N35), .B(N494), .Y(N678) );
  AND2X1 gate47 ( .A(N35), .B(N511), .Y(N681) );
  AND2X1 gate48 ( .A(N35), .B(N528), .Y(N684) );
  AND2X1 gate49 ( .A(N52), .B(N273), .Y(N687) );
  AND2X1 gate50 ( .A(N52), .B(N290), .Y(N690) );
  AND2X1 gate51 ( .A(N52), .B(N307), .Y(N693) );
  AND2X1 gate52 ( .A(N52), .B(N324), .Y(N696) );
  AND2X1 gate53 ( .A(N52), .B(N341), .Y(N699) );
  AND2X1 gate54 ( .A(N52), .B(N358), .Y(N702) );
  AND2X1 gate55 ( .A(N52), .B(N375), .Y(N705) );
  AND2X1 gate56 ( .A(N52), .B(N392), .Y(N708) );
  AND2X1 gate57 ( .A(N52), .B(N409), .Y(N711) );
  AND2X1 gate58 ( .A(N52), .B(N426), .Y(N714) );
  AND2X1 gate59 ( .A(N52), .B(N443), .Y(N717) );
  AND2X1 gate60 ( .A(N52), .B(N460), .Y(N720) );
  AND2X1 gate61 ( .A(N52), .B(N477), .Y(N723) );
  AND2X1 gate62 ( .A(N52), .B(N494), .Y(N726) );
  AND2X1 gate63 ( .A(N52), .B(N511), .Y(N729) );
  AND2X1 gate64 ( .A(N52), .B(N528), .Y(N732) );
  AND2X1 gate65 ( .A(N69), .B(N273), .Y(N735) );
  AND2X1 gate66 ( .A(N69), .B(N290), .Y(N738) );
  AND2X1 gate67 ( .A(N69), .B(N307), .Y(N741) );
  AND2X1 gate68 ( .A(N69), .B(N324), .Y(N744) );
  AND2X1 gate69 ( .A(N69), .B(N341), .Y(N747) );
  AND2X1 gate70 ( .A(N69), .B(N358), .Y(N750) );
  AND2X1 gate71 ( .A(N69), .B(N375), .Y(N753) );
  AND2X1 gate72 ( .A(N69), .B(N392), .Y(N756) );
  AND2X1 gate73 ( .A(N69), .B(N409), .Y(N759) );
  AND2X1 gate74 ( .A(N69), .B(N426), .Y(N762) );
  AND2X1 gate75 ( .A(N69), .B(N443), .Y(N765) );
  AND2X1 gate76 ( .A(N69), .B(N460), .Y(N768) );
  AND2X1 gate77 ( .A(N69), .B(N477), .Y(N771) );
  AND2X1 gate78 ( .A(N69), .B(N494), .Y(N774) );
  AND2X1 gate79 ( .A(N69), .B(N511), .Y(N777) );
  AND2X1 gate80 ( .A(N69), .B(N528), .Y(N780) );
  AND2X1 gate81 ( .A(N86), .B(N273), .Y(N783) );
  AND2X1 gate82 ( .A(N86), .B(N290), .Y(N786) );
  AND2X1 gate83 ( .A(N86), .B(N307), .Y(N789) );
  AND2X1 gate84 ( .A(N86), .B(N324), .Y(N792) );
  AND2X1 gate85 ( .A(N86), .B(N341), .Y(N795) );
  AND2X1 gate86 ( .A(N86), .B(N358), .Y(N798) );
  AND2X1 gate87 ( .A(N86), .B(N375), .Y(N801) );
  AND2X1 gate88 ( .A(N86), .B(N392), .Y(N804) );
  AND2X1 gate89 ( .A(N86), .B(N409), .Y(N807) );
  AND2X1 gate90 ( .A(N86), .B(N426), .Y(N810) );
  AND2X1 gate91 ( .A(N86), .B(N443), .Y(N813) );
  AND2X1 gate92 ( .A(N86), .B(N460), .Y(N816) );
  AND2X1 gate93 ( .A(N86), .B(N477), .Y(N819) );
  AND2X1 gate94 ( .A(N86), .B(N494), .Y(N822) );
  AND2X1 gate95 ( .A(N86), .B(N511), .Y(N825) );
  AND2X1 gate96 ( .A(N86), .B(N528), .Y(N828) );
  AND2X1 gate97 ( .A(N103), .B(N273), .Y(N831) );
  AND2X1 gate98 ( .A(N103), .B(N290), .Y(N834) );
  AND2X1 gate99 ( .A(N103), .B(N307), .Y(N837) );
  AND2X1 gate100 ( .A(N103), .B(N324), .Y(N840) );
  AND2X1 gate101 ( .A(N103), .B(N341), .Y(N843) );
  AND2X1 gate102 ( .A(N103), .B(N358), .Y(N846) );
  AND2X1 gate103 ( .A(N103), .B(N375), .Y(N849) );
  AND2X1 gate104 ( .A(N103), .B(N392), .Y(N852) );
  AND2X1 gate105 ( .A(N103), .B(N409), .Y(N855) );
  AND2X1 gate106 ( .A(N103), .B(N426), .Y(N858) );
  AND2X1 gate107 ( .A(N103), .B(N443), .Y(N861) );
  AND2X1 gate108 ( .A(N103), .B(N460), .Y(N864) );
  AND2X1 gate109 ( .A(N103), .B(N477), .Y(N867) );
  AND2X1 gate110 ( .A(N103), .B(N494), .Y(N870) );
  AND2X1 gate111 ( .A(N103), .B(N511), .Y(N873) );
  AND2X1 gate112 ( .A(N103), .B(N528), .Y(N876) );
  AND2X1 gate113 ( .A(N120), .B(N273), .Y(N879) );
  AND2X1 gate114 ( .A(N120), .B(N290), .Y(N882) );
  AND2X1 gate115 ( .A(N120), .B(N307), .Y(N885) );
  AND2X1 gate116 ( .A(N120), .B(N324), .Y(N888) );
  AND2X1 gate117 ( .A(N120), .B(N341), .Y(N891) );
  AND2X1 gate118 ( .A(N120), .B(N358), .Y(N894) );
  AND2X1 gate119 ( .A(N120), .B(N375), .Y(N897) );
  AND2X1 gate120 ( .A(N120), .B(N392), .Y(N900) );
  AND2X1 gate121 ( .A(N120), .B(N409), .Y(N903) );
  AND2X1 gate122 ( .A(N120), .B(N426), .Y(N906) );
  AND2X1 gate123 ( .A(N120), .B(N443), .Y(N909) );
  AND2X1 gate124 ( .A(N120), .B(N460), .Y(N912) );
  AND2X1 gate125 ( .A(N120), .B(N477), .Y(N915) );
  AND2X1 gate126 ( .A(N120), .B(N494), .Y(N918) );
  AND2X1 gate127 ( .A(N120), .B(N511), .Y(N921) );
  AND2X1 gate128 ( .A(N120), .B(N528), .Y(N924) );
  AND2X1 gate129 ( .A(N137), .B(N273), .Y(N927) );
  AND2X1 gate130 ( .A(N137), .B(N290), .Y(N930) );
  AND2X1 gate131 ( .A(N137), .B(N307), .Y(N933) );
  AND2X1 gate132 ( .A(N137), .B(N324), .Y(N936) );
  AND2X1 gate133 ( .A(N137), .B(N341), .Y(N939) );
  AND2X1 gate134 ( .A(N137), .B(N358), .Y(N942) );
  AND2X1 gate135 ( .A(N137), .B(N375), .Y(N945) );
  AND2X1 gate136 ( .A(N137), .B(N392), .Y(N948) );
  AND2X1 gate137 ( .A(N137), .B(N409), .Y(N951) );
  AND2X1 gate138 ( .A(N137), .B(N426), .Y(N954) );
  AND2X1 gate139 ( .A(N137), .B(N443), .Y(N957) );
  AND2X1 gate140 ( .A(N137), .B(N460), .Y(N960) );
  AND2X1 gate141 ( .A(N137), .B(N477), .Y(N963) );
  AND2X1 gate142 ( .A(N137), .B(N494), .Y(N966) );
  AND2X1 gate143 ( .A(N137), .B(N511), .Y(N969) );
  AND2X1 gate144 ( .A(N137), .B(N528), .Y(N972) );
  AND2X1 gate145 ( .A(N154), .B(N273), .Y(N975) );
  AND2X1 gate146 ( .A(N154), .B(N290), .Y(N978) );
  AND2X1 gate147 ( .A(N154), .B(N307), .Y(N981) );
  AND2X1 gate148 ( .A(N154), .B(N324), .Y(N984) );
  AND2X1 gate149 ( .A(N154), .B(N341), .Y(N987) );
  AND2X1 gate150 ( .A(N154), .B(N358), .Y(N990) );
  AND2X1 gate151 ( .A(N154), .B(N375), .Y(N993) );
  AND2X1 gate152 ( .A(N154), .B(N392), .Y(N996) );
  AND2X1 gate153 ( .A(N154), .B(N409), .Y(N999) );
  AND2X1 gate154 ( .A(N154), .B(N426), .Y(N1002) );
  AND2X1 gate155 ( .A(N154), .B(N443), .Y(N1005) );
  AND2X1 gate156 ( .A(N154), .B(N460), .Y(N1008) );
  AND2X1 gate157 ( .A(N154), .B(N477), .Y(N1011) );
  AND2X1 gate158 ( .A(N154), .B(N494), .Y(N1014) );
  AND2X1 gate159 ( .A(N154), .B(N511), .Y(N1017) );
  AND2X1 gate160 ( .A(N154), .B(N528), .Y(N1020) );
  AND2X1 gate161 ( .A(N171), .B(N273), .Y(N1023) );
  AND2X1 gate162 ( .A(N171), .B(N290), .Y(N1026) );
  AND2X1 gate163 ( .A(N171), .B(N307), .Y(N1029) );
  AND2X1 gate164 ( .A(N171), .B(N324), .Y(N1032) );
  AND2X1 gate165 ( .A(N171), .B(N341), .Y(N1035) );
  AND2X1 gate166 ( .A(N171), .B(N358), .Y(N1038) );
  AND2X1 gate167 ( .A(N171), .B(N375), .Y(N1041) );
  AND2X1 gate168 ( .A(N171), .B(N392), .Y(N1044) );
  AND2X1 gate169 ( .A(N171), .B(N409), .Y(N1047) );
  AND2X1 gate170 ( .A(N171), .B(N426), .Y(N1050) );
  AND2X1 gate171 ( .A(N171), .B(N443), .Y(N1053) );
  AND2X1 gate172 ( .A(N171), .B(N460), .Y(N1056) );
  AND2X1 gate173 ( .A(N171), .B(N477), .Y(N1059) );
  AND2X1 gate174 ( .A(N171), .B(N494), .Y(N1062) );
  AND2X1 gate175 ( .A(N171), .B(N511), .Y(N1065) );
  AND2X1 gate176 ( .A(N171), .B(N528), .Y(N1068) );
  AND2X1 gate177 ( .A(N188), .B(N273), .Y(N1071) );
  AND2X1 gate178 ( .A(N188), .B(N290), .Y(N1074) );
  AND2X1 gate179 ( .A(N188), .B(N307), .Y(N1077) );
  AND2X1 gate180 ( .A(N188), .B(N324), .Y(N1080) );
  AND2X1 gate181 ( .A(N188), .B(N341), .Y(N1083) );
  AND2X1 gate182 ( .A(N188), .B(N358), .Y(N1086) );
  AND2X1 gate183 ( .A(N188), .B(N375), .Y(N1089) );
  AND2X1 gate184 ( .A(N188), .B(N392), .Y(N1092) );
  AND2X1 gate185 ( .A(N188), .B(N409), .Y(N1095) );
  AND2X1 gate186 ( .A(N188), .B(N426), .Y(N1098) );
  AND2X1 gate187 ( .A(N188), .B(N443), .Y(N1101) );
  AND2X1 gate188 ( .A(N188), .B(N460), .Y(N1104) );
  AND2X1 gate189 ( .A(N188), .B(N477), .Y(N1107) );
  AND2X1 gate190 ( .A(N188), .B(N494), .Y(N1110) );
  AND2X1 gate191 ( .A(N188), .B(N511), .Y(N1113) );
  AND2X1 gate192 ( .A(N188), .B(N528), .Y(N1116) );
  AND2X1 gate193 ( .A(N205), .B(N273), .Y(N1119) );
  AND2X1 gate194 ( .A(N205), .B(N290), .Y(N1122) );
  AND2X1 gate195 ( .A(N205), .B(N307), .Y(N1125) );
  AND2X1 gate196 ( .A(N205), .B(N324), .Y(N1128) );
  AND2X1 gate197 ( .A(N205), .B(N341), .Y(N1131) );
  AND2X1 gate198 ( .A(N205), .B(N358), .Y(N1134) );
  AND2X1 gate199 ( .A(N205), .B(N375), .Y(N1137) );
  AND2X1 gate200 ( .A(N205), .B(N392), .Y(N1140) );
  AND2X1 gate201 ( .A(N205), .B(N409), .Y(N1143) );
  AND2X1 gate202 ( .A(N205), .B(N426), .Y(N1146) );
  AND2X1 gate203 ( .A(N205), .B(N443), .Y(N1149) );
  AND2X1 gate204 ( .A(N205), .B(N460), .Y(N1152) );
  AND2X1 gate205 ( .A(N205), .B(N477), .Y(N1155) );
  AND2X1 gate206 ( .A(N205), .B(N494), .Y(N1158) );
  AND2X1 gate207 ( .A(N205), .B(N511), .Y(N1161) );
  AND2X1 gate208 ( .A(N205), .B(N528), .Y(N1164) );
  AND2X1 gate209 ( .A(N222), .B(N273), .Y(N1167) );
  AND2X1 gate210 ( .A(N222), .B(N290), .Y(N1170) );
  AND2X1 gate211 ( .A(N222), .B(N307), .Y(N1173) );
  AND2X1 gate212 ( .A(N222), .B(N324), .Y(N1176) );
  AND2X1 gate213 ( .A(N222), .B(N341), .Y(N1179) );
  AND2X1 gate214 ( .A(N222), .B(N358), .Y(N1182) );
  AND2X1 gate215 ( .A(N222), .B(N375), .Y(N1185) );
  AND2X1 gate216 ( .A(N222), .B(N392), .Y(N1188) );
  AND2X1 gate217 ( .A(N222), .B(N409), .Y(N1191) );
  AND2X1 gate218 ( .A(N222), .B(N426), .Y(N1194) );
  AND2X1 gate219 ( .A(N222), .B(N443), .Y(N1197) );
  AND2X1 gate220 ( .A(N222), .B(N460), .Y(N1200) );
  AND2X1 gate221 ( .A(N222), .B(N477), .Y(N1203) );
  AND2X1 gate222 ( .A(N222), .B(N494), .Y(N1206) );
  AND2X1 gate223 ( .A(N222), .B(N511), .Y(N1209) );
  AND2X1 gate224 ( .A(N222), .B(N528), .Y(N1212) );
  AND2X1 gate225 ( .A(N239), .B(N273), .Y(N1215) );
  AND2X1 gate226 ( .A(N239), .B(N290), .Y(N1218) );
  AND2X1 gate227 ( .A(N239), .B(N307), .Y(N1221) );
  AND2X1 gate228 ( .A(N239), .B(N324), .Y(N1224) );
  AND2X1 gate229 ( .A(N239), .B(N341), .Y(N1227) );
  AND2X1 gate230 ( .A(N239), .B(N358), .Y(N1230) );
  AND2X1 gate231 ( .A(N239), .B(N375), .Y(N1233) );
  AND2X1 gate232 ( .A(N239), .B(N392), .Y(N1236) );
  AND2X1 gate233 ( .A(N239), .B(N409), .Y(N1239) );
  AND2X1 gate234 ( .A(N239), .B(N426), .Y(N1242) );
  AND2X1 gate235 ( .A(N239), .B(N443), .Y(N1245) );
  AND2X1 gate236 ( .A(N239), .B(N460), .Y(N1248) );
  AND2X1 gate237 ( .A(N239), .B(N477), .Y(N1251) );
  AND2X1 gate238 ( .A(N239), .B(N494), .Y(N1254) );
  AND2X1 gate239 ( .A(N239), .B(N511), .Y(N1257) );
  AND2X1 gate240 ( .A(N239), .B(N528), .Y(N1260) );
  AND2X1 gate241 ( .A(N256), .B(N273), .Y(N1263) );
  AND2X1 gate242 ( .A(N256), .B(N290), .Y(N1266) );
  AND2X1 gate243 ( .A(N256), .B(N307), .Y(N1269) );
  AND2X1 gate244 ( .A(N256), .B(N324), .Y(N1272) );
  AND2X1 gate245 ( .A(N256), .B(N341), .Y(N1275) );
  AND2X1 gate246 ( .A(N256), .B(N358), .Y(N1278) );
  AND2X1 gate247 ( .A(N256), .B(N375), .Y(N1281) );
  AND2X1 gate248 ( .A(N256), .B(N392), .Y(N1284) );
  AND2X1 gate249 ( .A(N256), .B(N409), .Y(N1287) );
  AND2X1 gate250 ( .A(N256), .B(N426), .Y(N1290) );
  AND2X1 gate251 ( .A(N256), .B(N443), .Y(N1293) );
  AND2X1 gate252 ( .A(N256), .B(N460), .Y(N1296) );
  AND2X1 gate253 ( .A(N256), .B(N477), .Y(N1299) );
  AND2X1 gate254 ( .A(N256), .B(N494), .Y(N1302) );
  AND2X1 gate255 ( .A(N256), .B(N511), .Y(N1305) );
  AND2X1 gate256 ( .A(N256), .B(N528), .Y(N1308) );
  INVX1 gate257 ( .A(N591), .Y(N1311) );
  INVX1 gate258 ( .A(N639), .Y(N1315) );
  INVX1 gate259 ( .A(N687), .Y(N1319) );
  INVX1 gate260 ( .A(N735), .Y(N1323) );
  INVX1 gate261 ( .A(N783), .Y(N1327) );
  INVX1 gate262 ( .A(N831), .Y(N1331) );
  INVX1 gate263 ( .A(N879), .Y(N1335) );
  INVX1 gate264 ( .A(N927), .Y(N1339) );
  INVX1 gate265 ( .A(N975), .Y(N1343) );
  INVX1 gate266 ( .A(N1023), .Y(N1347) );
  INVX1 gate267 ( .A(N1071), .Y(N1351) );
  INVX1 gate268 ( .A(N1119), .Y(N1355) );
  INVX1 gate269 ( .A(N1167), .Y(N1359) );
  INVX1 gate270 ( .A(N1215), .Y(N1363) );
  INVX1 gate271 ( .A(N1263), .Y(N1367) );
  NOR2X1 gate272 ( .A(N591), .B(N1311), .Y(N1371) );
  INVX1 gate273 ( .A(N1311), .Y(N1372) );
  NOR2X1 gate274 ( .A(N639), .B(N1315), .Y(N1373) );
  INVX1 gate275 ( .A(N1315), .Y(N1374) );
  NOR2X1 gate276 ( .A(N687), .B(N1319), .Y(N1375) );
  INVX1 gate277 ( .A(N1319), .Y(N1376) );
  NOR2X1 gate278 ( .A(N735), .B(N1323), .Y(N1377) );
  INVX1 gate279 ( .A(N1323), .Y(N1378) );
  NOR2X1 gate280 ( .A(N783), .B(N1327), .Y(N1379) );
  INVX1 gate281 ( .A(N1327), .Y(N1380) );
  NOR2X1 gate282 ( .A(N831), .B(N1331), .Y(N1381) );
  INVX1 gate283 ( .A(N1331), .Y(N1382) );
  NOR2X1 gate284 ( .A(N879), .B(N1335), .Y(N1383) );
  INVX1 gate285 ( .A(N1335), .Y(N1384) );
  NOR2X1 gate286 ( .A(N927), .B(N1339), .Y(N1385) );
  INVX1 gate287 ( .A(N1339), .Y(N1386) );
  NOR2X1 gate288 ( .A(N975), .B(N1343), .Y(N1387) );
  INVX1 gate289 ( .A(N1343), .Y(N1388) );
  NOR2X1 gate290 ( .A(N1023), .B(N1347), .Y(N1389) );
  INVX1 gate291 ( .A(N1347), .Y(N1390) );
  NOR2X1 gate292 ( .A(N1071), .B(N1351), .Y(N1391) );
  INVX1 gate293 ( .A(N1351), .Y(N1392) );
  NOR2X1 gate294 ( .A(N1119), .B(N1355), .Y(N1393) );
  INVX1 gate295 ( .A(N1355), .Y(N1394) );
  NOR2X1 gate296 ( .A(N1167), .B(N1359), .Y(N1395) );
  INVX1 gate297 ( .A(N1359), .Y(N1396) );
  NOR2X1 gate298 ( .A(N1215), .B(N1363), .Y(N1397) );
  INVX1 gate299 ( .A(N1363), .Y(N1398) );
  NOR2X1 gate300 ( .A(N1263), .B(N1367), .Y(N1399) );
  INVX1 gate301 ( .A(N1367), .Y(N1400) );
  NOR2X1 gate302 ( .A(N1371), .B(N1372), .Y(N1401) );
  NOR2X1 gate303 ( .A(N1373), .B(N1374), .Y(N1404) );
  NOR2X1 gate304 ( .A(N1375), .B(N1376), .Y(N1407) );
  NOR2X1 gate305 ( .A(N1377), .B(N1378), .Y(N1410) );
  NOR2X1 gate306 ( .A(N1379), .B(N1380), .Y(N1413) );
  NOR2X1 gate307 ( .A(N1381), .B(N1382), .Y(N1416) );
  NOR2X1 gate308 ( .A(N1383), .B(N1384), .Y(N1419) );
  NOR2X1 gate309 ( .A(N1385), .B(N1386), .Y(N1422) );
  NOR2X1 gate310 ( .A(N1387), .B(N1388), .Y(N1425) );
  NOR2X1 gate311 ( .A(N1389), .B(N1390), .Y(N1428) );
  NOR2X1 gate312 ( .A(N1391), .B(N1392), .Y(N1431) );
  NOR2X1 gate313 ( .A(N1393), .B(N1394), .Y(N1434) );
  NOR2X1 gate314 ( .A(N1395), .B(N1396), .Y(N1437) );
  NOR2X1 gate315 ( .A(N1397), .B(N1398), .Y(N1440) );
  NOR2X1 gate316 ( .A(N1399), .B(N1400), .Y(N1443) );
  NOR2X1 gate317 ( .A(N1401), .B(N546), .Y(N1446) );
  NOR2X1 gate318 ( .A(N1404), .B(N594), .Y(N1450) );
  NOR2X1 gate319 ( .A(N1407), .B(N642), .Y(N1454) );
  NOR2X1 gate320 ( .A(N1410), .B(N690), .Y(N1458) );
  NOR2X1 gate321 ( .A(N1413), .B(N738), .Y(N1462) );
  NOR2X1 gate322 ( .A(N1416), .B(N786), .Y(N1466) );
  NOR2X1 gate323 ( .A(N1419), .B(N834), .Y(N1470) );
  NOR2X1 gate324 ( .A(N1422), .B(N882), .Y(N1474) );
  NOR2X1 gate325 ( .A(N1425), .B(N930), .Y(N1478) );
  NOR2X1 gate326 ( .A(N1428), .B(N978), .Y(N1482) );
  NOR2X1 gate327 ( .A(N1431), .B(N1026), .Y(N1486) );
  NOR2X1 gate328 ( .A(N1434), .B(N1074), .Y(N1490) );
  NOR2X1 gate329 ( .A(N1437), .B(N1122), .Y(N1494) );
  NOR2X1 gate330 ( .A(N1440), .B(N1170), .Y(N1498) );
  NOR2X1 gate331 ( .A(N1443), .B(N1218), .Y(N1502) );
  NOR2X1 gate332 ( .A(N1401), .B(N1446), .Y(N1506) );
  NOR2X1 gate333 ( .A(N1446), .B(N546), .Y(N1507) );
  NOR2X1 gate334 ( .A(N1311), .B(N1446), .Y(N1508) );
  NOR2X1 gate335 ( .A(N1404), .B(N1450), .Y(N1511) );
  NOR2X1 gate336 ( .A(N1450), .B(N594), .Y(N1512) );
  NOR2X1 gate337 ( .A(N1315), .B(N1450), .Y(N1513) );
  NOR2X1 gate338 ( .A(N1407), .B(N1454), .Y(N1516) );
  NOR2X1 gate339 ( .A(N1454), .B(N642), .Y(N1517) );
  NOR2X1 gate340 ( .A(N1319), .B(N1454), .Y(N1518) );
  NOR2X1 gate341 ( .A(N1410), .B(N1458), .Y(N1521) );
  NOR2X1 gate342 ( .A(N1458), .B(N690), .Y(N1522) );
  NOR2X1 gate343 ( .A(N1323), .B(N1458), .Y(N1523) );
  NOR2X1 gate344 ( .A(N1413), .B(N1462), .Y(N1526) );
  NOR2X1 gate345 ( .A(N1462), .B(N738), .Y(N1527) );
  NOR2X1 gate346 ( .A(N1327), .B(N1462), .Y(N1528) );
  NOR2X1 gate347 ( .A(N1416), .B(N1466), .Y(N1531) );
  NOR2X1 gate348 ( .A(N1466), .B(N786), .Y(N1532) );
  NOR2X1 gate349 ( .A(N1331), .B(N1466), .Y(N1533) );
  NOR2X1 gate350 ( .A(N1419), .B(N1470), .Y(N1536) );
  NOR2X1 gate351 ( .A(N1470), .B(N834), .Y(N1537) );
  NOR2X1 gate352 ( .A(N1335), .B(N1470), .Y(N1538) );
  NOR2X1 gate353 ( .A(N1422), .B(N1474), .Y(N1541) );
  NOR2X1 gate354 ( .A(N1474), .B(N882), .Y(N1542) );
  NOR2X1 gate355 ( .A(N1339), .B(N1474), .Y(N1543) );
  NOR2X1 gate356 ( .A(N1425), .B(N1478), .Y(N1546) );
  NOR2X1 gate357 ( .A(N1478), .B(N930), .Y(N1547) );
  NOR2X1 gate358 ( .A(N1343), .B(N1478), .Y(N1548) );
  NOR2X1 gate359 ( .A(N1428), .B(N1482), .Y(N1551) );
  NOR2X1 gate360 ( .A(N1482), .B(N978), .Y(N1552) );
  NOR2X1 gate361 ( .A(N1347), .B(N1482), .Y(N1553) );
  NOR2X1 gate362 ( .A(N1431), .B(N1486), .Y(N1556) );
  NOR2X1 gate363 ( .A(N1486), .B(N1026), .Y(N1557) );
  NOR2X1 gate364 ( .A(N1351), .B(N1486), .Y(N1558) );
  NOR2X1 gate365 ( .A(N1434), .B(N1490), .Y(N1561) );
  NOR2X1 gate366 ( .A(N1490), .B(N1074), .Y(N1562) );
  NOR2X1 gate367 ( .A(N1355), .B(N1490), .Y(N1563) );
  NOR2X1 gate368 ( .A(N1437), .B(N1494), .Y(N1566) );
  NOR2X1 gate369 ( .A(N1494), .B(N1122), .Y(N1567) );
  NOR2X1 gate370 ( .A(N1359), .B(N1494), .Y(N1568) );
  NOR2X1 gate371 ( .A(N1440), .B(N1498), .Y(N1571) );
  NOR2X1 gate372 ( .A(N1498), .B(N1170), .Y(N1572) );
  NOR2X1 gate373 ( .A(N1363), .B(N1498), .Y(N1573) );
  NOR2X1 gate374 ( .A(N1443), .B(N1502), .Y(N1576) );
  NOR2X1 gate375 ( .A(N1502), .B(N1218), .Y(N1577) );
  NOR2X1 gate376 ( .A(N1367), .B(N1502), .Y(N1578) );
  NOR2X1 gate377 ( .A(N1506), .B(N1507), .Y(N1581) );
  NOR2X1 gate378 ( .A(N1511), .B(N1512), .Y(N1582) );
  NOR2X1 gate379 ( .A(N1516), .B(N1517), .Y(N1585) );
  NOR2X1 gate380 ( .A(N1521), .B(N1522), .Y(N1588) );
  NOR2X1 gate381 ( .A(N1526), .B(N1527), .Y(N1591) );
  NOR2X1 gate382 ( .A(N1531), .B(N1532), .Y(N1594) );
  NOR2X1 gate383 ( .A(N1536), .B(N1537), .Y(N1597) );
  NOR2X1 gate384 ( .A(N1541), .B(N1542), .Y(N1600) );
  NOR2X1 gate385 ( .A(N1546), .B(N1547), .Y(N1603) );
  NOR2X1 gate386 ( .A(N1551), .B(N1552), .Y(N1606) );
  NOR2X1 gate387 ( .A(N1556), .B(N1557), .Y(N1609) );
  NOR2X1 gate388 ( .A(N1561), .B(N1562), .Y(N1612) );
  NOR2X1 gate389 ( .A(N1566), .B(N1567), .Y(N1615) );
  NOR2X1 gate390 ( .A(N1571), .B(N1572), .Y(N1618) );
  NOR2X1 gate391 ( .A(N1576), .B(N1577), .Y(N1621) );
  NOR2X1 gate392 ( .A(N1266), .B(N1578), .Y(N1624) );
  NOR2X1 gate393 ( .A(N1582), .B(N1508), .Y(N1628) );
  NOR2X1 gate394 ( .A(N1585), .B(N1513), .Y(N1632) );
  NOR2X1 gate395 ( .A(N1588), .B(N1518), .Y(N1636) );
  NOR2X1 gate396 ( .A(N1591), .B(N1523), .Y(N1640) );
  NOR2X1 gate397 ( .A(N1594), .B(N1528), .Y(N1644) );
  NOR2X1 gate398 ( .A(N1597), .B(N1533), .Y(N1648) );
  NOR2X1 gate399 ( .A(N1600), .B(N1538), .Y(N1652) );
  NOR2X1 gate400 ( .A(N1603), .B(N1543), .Y(N1656) );
  NOR2X1 gate401 ( .A(N1606), .B(N1548), .Y(N1660) );
  NOR2X1 gate402 ( .A(N1609), .B(N1553), .Y(N1664) );
  NOR2X1 gate403 ( .A(N1612), .B(N1558), .Y(N1668) );
  NOR2X1 gate404 ( .A(N1615), .B(N1563), .Y(N1672) );
  NOR2X1 gate405 ( .A(N1618), .B(N1568), .Y(N1676) );
  NOR2X1 gate406 ( .A(N1621), .B(N1573), .Y(N1680) );
  NOR2X1 gate407 ( .A(N1266), .B(N1624), .Y(N1684) );
  NOR2X1 gate408 ( .A(N1624), .B(N1578), .Y(N1685) );
  NOR2X1 gate409 ( .A(N1582), .B(N1628), .Y(N1686) );
  NOR2X1 gate410 ( .A(N1628), .B(N1508), .Y(N1687) );
  NOR2X1 gate411 ( .A(N1585), .B(N1632), .Y(N1688) );
  NOR2X1 gate412 ( .A(N1632), .B(N1513), .Y(N1689) );
  NOR2X1 gate413 ( .A(N1588), .B(N1636), .Y(N1690) );
  NOR2X1 gate414 ( .A(N1636), .B(N1518), .Y(N1691) );
  NOR2X1 gate415 ( .A(N1591), .B(N1640), .Y(N1692) );
  NOR2X1 gate416 ( .A(N1640), .B(N1523), .Y(N1693) );
  NOR2X1 gate417 ( .A(N1594), .B(N1644), .Y(N1694) );
  NOR2X1 gate418 ( .A(N1644), .B(N1528), .Y(N1695) );
  NOR2X1 gate419 ( .A(N1597), .B(N1648), .Y(N1696) );
  NOR2X1 gate420 ( .A(N1648), .B(N1533), .Y(N1697) );
  NOR2X1 gate421 ( .A(N1600), .B(N1652), .Y(N1698) );
  NOR2X1 gate422 ( .A(N1652), .B(N1538), .Y(N1699) );
  NOR2X1 gate423 ( .A(N1603), .B(N1656), .Y(N1700) );
  NOR2X1 gate424 ( .A(N1656), .B(N1543), .Y(N1701) );
  NOR2X1 gate425 ( .A(N1606), .B(N1660), .Y(N1702) );
  NOR2X1 gate426 ( .A(N1660), .B(N1548), .Y(N1703) );
  NOR2X1 gate427 ( .A(N1609), .B(N1664), .Y(N1704) );
  NOR2X1 gate428 ( .A(N1664), .B(N1553), .Y(N1705) );
  NOR2X1 gate429 ( .A(N1612), .B(N1668), .Y(N1706) );
  NOR2X1 gate430 ( .A(N1668), .B(N1558), .Y(N1707) );
  NOR2X1 gate431 ( .A(N1615), .B(N1672), .Y(N1708) );
  NOR2X1 gate432 ( .A(N1672), .B(N1563), .Y(N1709) );
  NOR2X1 gate433 ( .A(N1618), .B(N1676), .Y(N1710) );
  NOR2X1 gate434 ( .A(N1676), .B(N1568), .Y(N1711) );
  NOR2X1 gate435 ( .A(N1621), .B(N1680), .Y(N1712) );
  NOR2X1 gate436 ( .A(N1680), .B(N1573), .Y(N1713) );
  NOR2X1 gate437 ( .A(N1684), .B(N1685), .Y(N1714) );
  NOR2X1 gate438 ( .A(N1686), .B(N1687), .Y(N1717) );
  NOR2X1 gate439 ( .A(N1688), .B(N1689), .Y(N1720) );
  NOR2X1 gate440 ( .A(N1690), .B(N1691), .Y(N1723) );
  NOR2X1 gate441 ( .A(N1692), .B(N1693), .Y(N1726) );
  NOR2X1 gate442 ( .A(N1694), .B(N1695), .Y(N1729) );
  NOR2X1 gate443 ( .A(N1696), .B(N1697), .Y(N1732) );
  NOR2X1 gate444 ( .A(N1698), .B(N1699), .Y(N1735) );
  NOR2X1 gate445 ( .A(N1700), .B(N1701), .Y(N1738) );
  NOR2X1 gate446 ( .A(N1702), .B(N1703), .Y(N1741) );
  NOR2X1 gate447 ( .A(N1704), .B(N1705), .Y(N1744) );
  NOR2X1 gate448 ( .A(N1706), .B(N1707), .Y(N1747) );
  NOR2X1 gate449 ( .A(N1708), .B(N1709), .Y(N1750) );
  NOR2X1 gate450 ( .A(N1710), .B(N1711), .Y(N1753) );
  NOR2X1 gate451 ( .A(N1712), .B(N1713), .Y(N1756) );
  NOR2X1 gate452 ( .A(N1714), .B(N1221), .Y(N1759) );
  NOR2X1 gate453 ( .A(N1717), .B(N549), .Y(N1763) );
  NOR2X1 gate454 ( .A(N1720), .B(N597), .Y(N1767) );
  NOR2X1 gate455 ( .A(N1723), .B(N645), .Y(N1771) );
  NOR2X1 gate456 ( .A(N1726), .B(N693), .Y(N1775) );
  NOR2X1 gate457 ( .A(N1729), .B(N741), .Y(N1779) );
  NOR2X1 gate458 ( .A(N1732), .B(N789), .Y(N1783) );
  NOR2X1 gate459 ( .A(N1735), .B(N837), .Y(N1787) );
  NOR2X1 gate460 ( .A(N1738), .B(N885), .Y(N1791) );
  NOR2X1 gate461 ( .A(N1741), .B(N933), .Y(N1795) );
  NOR2X1 gate462 ( .A(N1744), .B(N981), .Y(N1799) );
  NOR2X1 gate463 ( .A(N1747), .B(N1029), .Y(N1803) );
  NOR2X1 gate464 ( .A(N1750), .B(N1077), .Y(N1807) );
  NOR2X1 gate465 ( .A(N1753), .B(N1125), .Y(N1811) );
  NOR2X1 gate466 ( .A(N1756), .B(N1173), .Y(N1815) );
  NOR2X1 gate467 ( .A(N1714), .B(N1759), .Y(N1819) );
  NOR2X1 gate468 ( .A(N1759), .B(N1221), .Y(N1820) );
  NOR2X1 gate469 ( .A(N1624), .B(N1759), .Y(N1821) );
  NOR2X1 gate470 ( .A(N1717), .B(N1763), .Y(N1824) );
  NOR2X1 gate471 ( .A(N1763), .B(N549), .Y(N1825) );
  NOR2X1 gate472 ( .A(N1628), .B(N1763), .Y(N1826) );
  NOR2X1 gate473 ( .A(N1720), .B(N1767), .Y(N1829) );
  NOR2X1 gate474 ( .A(N1767), .B(N597), .Y(N1830) );
  NOR2X1 gate475 ( .A(N1632), .B(N1767), .Y(N1831) );
  NOR2X1 gate476 ( .A(N1723), .B(N1771), .Y(N1834) );
  NOR2X1 gate477 ( .A(N1771), .B(N645), .Y(N1835) );
  NOR2X1 gate478 ( .A(N1636), .B(N1771), .Y(N1836) );
  NOR2X1 gate479 ( .A(N1726), .B(N1775), .Y(N1839) );
  NOR2X1 gate480 ( .A(N1775), .B(N693), .Y(N1840) );
  NOR2X1 gate481 ( .A(N1640), .B(N1775), .Y(N1841) );
  NOR2X1 gate482 ( .A(N1729), .B(N1779), .Y(N1844) );
  NOR2X1 gate483 ( .A(N1779), .B(N741), .Y(N1845) );
  NOR2X1 gate484 ( .A(N1644), .B(N1779), .Y(N1846) );
  NOR2X1 gate485 ( .A(N1732), .B(N1783), .Y(N1849) );
  NOR2X1 gate486 ( .A(N1783), .B(N789), .Y(N1850) );
  NOR2X1 gate487 ( .A(N1648), .B(N1783), .Y(N1851) );
  NOR2X1 gate488 ( .A(N1735), .B(N1787), .Y(N1854) );
  NOR2X1 gate489 ( .A(N1787), .B(N837), .Y(N1855) );
  NOR2X1 gate490 ( .A(N1652), .B(N1787), .Y(N1856) );
  NOR2X1 gate491 ( .A(N1738), .B(N1791), .Y(N1859) );
  NOR2X1 gate492 ( .A(N1791), .B(N885), .Y(N1860) );
  NOR2X1 gate493 ( .A(N1656), .B(N1791), .Y(N1861) );
  NOR2X1 gate494 ( .A(N1741), .B(N1795), .Y(N1864) );
  NOR2X1 gate495 ( .A(N1795), .B(N933), .Y(N1865) );
  NOR2X1 gate496 ( .A(N1660), .B(N1795), .Y(N1866) );
  NOR2X1 gate497 ( .A(N1744), .B(N1799), .Y(N1869) );
  NOR2X1 gate498 ( .A(N1799), .B(N981), .Y(N1870) );
  NOR2X1 gate499 ( .A(N1664), .B(N1799), .Y(N1871) );
  NOR2X1 gate500 ( .A(N1747), .B(N1803), .Y(N1874) );
  NOR2X1 gate501 ( .A(N1803), .B(N1029), .Y(N1875) );
  NOR2X1 gate502 ( .A(N1668), .B(N1803), .Y(N1876) );
  NOR2X1 gate503 ( .A(N1750), .B(N1807), .Y(N1879) );
  NOR2X1 gate504 ( .A(N1807), .B(N1077), .Y(N1880) );
  NOR2X1 gate505 ( .A(N1672), .B(N1807), .Y(N1881) );
  NOR2X1 gate506 ( .A(N1753), .B(N1811), .Y(N1884) );
  NOR2X1 gate507 ( .A(N1811), .B(N1125), .Y(N1885) );
  NOR2X1 gate508 ( .A(N1676), .B(N1811), .Y(N1886) );
  NOR2X1 gate509 ( .A(N1756), .B(N1815), .Y(N1889) );
  NOR2X1 gate510 ( .A(N1815), .B(N1173), .Y(N1890) );
  NOR2X1 gate511 ( .A(N1680), .B(N1815), .Y(N1891) );
  NOR2X1 gate512 ( .A(N1819), .B(N1820), .Y(N1894) );
  NOR2X1 gate513 ( .A(N1269), .B(N1821), .Y(N1897) );
  NOR2X1 gate514 ( .A(N1824), .B(N1825), .Y(N1901) );
  NOR2X1 gate515 ( .A(N1829), .B(N1830), .Y(N1902) );
  NOR2X1 gate516 ( .A(N1834), .B(N1835), .Y(N1905) );
  NOR2X1 gate517 ( .A(N1839), .B(N1840), .Y(N1908) );
  NOR2X1 gate518 ( .A(N1844), .B(N1845), .Y(N1911) );
  NOR2X1 gate519 ( .A(N1849), .B(N1850), .Y(N1914) );
  NOR2X1 gate520 ( .A(N1854), .B(N1855), .Y(N1917) );
  NOR2X1 gate521 ( .A(N1859), .B(N1860), .Y(N1920) );
  NOR2X1 gate522 ( .A(N1864), .B(N1865), .Y(N1923) );
  NOR2X1 gate523 ( .A(N1869), .B(N1870), .Y(N1926) );
  NOR2X1 gate524 ( .A(N1874), .B(N1875), .Y(N1929) );
  NOR2X1 gate525 ( .A(N1879), .B(N1880), .Y(N1932) );
  NOR2X1 gate526 ( .A(N1884), .B(N1885), .Y(N1935) );
  NOR2X1 gate527 ( .A(N1889), .B(N1890), .Y(N1938) );
  NOR2X1 gate528 ( .A(N1894), .B(N1891), .Y(N1941) );
  NOR2X1 gate529 ( .A(N1269), .B(N1897), .Y(N1945) );
  NOR2X1 gate530 ( .A(N1897), .B(N1821), .Y(N1946) );
  NOR2X1 gate531 ( .A(N1902), .B(N1826), .Y(N1947) );
  NOR2X1 gate532 ( .A(N1905), .B(N1831), .Y(N1951) );
  NOR2X1 gate533 ( .A(N1908), .B(N1836), .Y(N1955) );
  NOR2X1 gate534 ( .A(N1911), .B(N1841), .Y(N1959) );
  NOR2X1 gate535 ( .A(N1914), .B(N1846), .Y(N1963) );
  NOR2X1 gate536 ( .A(N1917), .B(N1851), .Y(N1967) );
  NOR2X1 gate537 ( .A(N1920), .B(N1856), .Y(N1971) );
  NOR2X1 gate538 ( .A(N1923), .B(N1861), .Y(N1975) );
  NOR2X1 gate539 ( .A(N1926), .B(N1866), .Y(N1979) );
  NOR2X1 gate540 ( .A(N1929), .B(N1871), .Y(N1983) );
  NOR2X1 gate541 ( .A(N1932), .B(N1876), .Y(N1987) );
  NOR2X1 gate542 ( .A(N1935), .B(N1881), .Y(N1991) );
  NOR2X1 gate543 ( .A(N1938), .B(N1886), .Y(N1995) );
  NOR2X1 gate544 ( .A(N1894), .B(N1941), .Y(N1999) );
  NOR2X1 gate545 ( .A(N1941), .B(N1891), .Y(N2000) );
  NOR2X1 gate546 ( .A(N1945), .B(N1946), .Y(N2001) );
  NOR2X1 gate547 ( .A(N1902), .B(N1947), .Y(N2004) );
  NOR2X1 gate548 ( .A(N1947), .B(N1826), .Y(N2005) );
  NOR2X1 gate549 ( .A(N1905), .B(N1951), .Y(N2006) );
  NOR2X1 gate550 ( .A(N1951), .B(N1831), .Y(N2007) );
  NOR2X1 gate551 ( .A(N1908), .B(N1955), .Y(N2008) );
  NOR2X1 gate552 ( .A(N1955), .B(N1836), .Y(N2009) );
  NOR2X1 gate553 ( .A(N1911), .B(N1959), .Y(N2010) );
  NOR2X1 gate554 ( .A(N1959), .B(N1841), .Y(N2011) );
  NOR2X1 gate555 ( .A(N1914), .B(N1963), .Y(N2012) );
  NOR2X1 gate556 ( .A(N1963), .B(N1846), .Y(N2013) );
  NOR2X1 gate557 ( .A(N1917), .B(N1967), .Y(N2014) );
  NOR2X1 gate558 ( .A(N1967), .B(N1851), .Y(N2015) );
  NOR2X1 gate559 ( .A(N1920), .B(N1971), .Y(N2016) );
  NOR2X1 gate560 ( .A(N1971), .B(N1856), .Y(N2017) );
  NOR2X1 gate561 ( .A(N1923), .B(N1975), .Y(N2018) );
  NOR2X1 gate562 ( .A(N1975), .B(N1861), .Y(N2019) );
  NOR2X1 gate563 ( .A(N1926), .B(N1979), .Y(N2020) );
  NOR2X1 gate564 ( .A(N1979), .B(N1866), .Y(N2021) );
  NOR2X1 gate565 ( .A(N1929), .B(N1983), .Y(N2022) );
  NOR2X1 gate566 ( .A(N1983), .B(N1871), .Y(N2023) );
  NOR2X1 gate567 ( .A(N1932), .B(N1987), .Y(N2024) );
  NOR2X1 gate568 ( .A(N1987), .B(N1876), .Y(N2025) );
  NOR2X1 gate569 ( .A(N1935), .B(N1991), .Y(N2026) );
  NOR2X1 gate570 ( .A(N1991), .B(N1881), .Y(N2027) );
  NOR2X1 gate571 ( .A(N1938), .B(N1995), .Y(N2028) );
  NOR2X1 gate572 ( .A(N1995), .B(N1886), .Y(N2029) );
  NOR2X1 gate573 ( .A(N1999), .B(N2000), .Y(N2030) );
  NOR2X1 gate574 ( .A(N2001), .B(N1224), .Y(N2033) );
  NOR2X1 gate575 ( .A(N2004), .B(N2005), .Y(N2037) );
  NOR2X1 gate576 ( .A(N2006), .B(N2007), .Y(N2040) );
  NOR2X1 gate577 ( .A(N2008), .B(N2009), .Y(N2043) );
  NOR2X1 gate578 ( .A(N2010), .B(N2011), .Y(N2046) );
  NOR2X1 gate579 ( .A(N2012), .B(N2013), .Y(N2049) );
  NOR2X1 gate580 ( .A(N2014), .B(N2015), .Y(N2052) );
  NOR2X1 gate581 ( .A(N2016), .B(N2017), .Y(N2055) );
  NOR2X1 gate582 ( .A(N2018), .B(N2019), .Y(N2058) );
  NOR2X1 gate583 ( .A(N2020), .B(N2021), .Y(N2061) );
  NOR2X1 gate584 ( .A(N2022), .B(N2023), .Y(N2064) );
  NOR2X1 gate585 ( .A(N2024), .B(N2025), .Y(N2067) );
  NOR2X1 gate586 ( .A(N2026), .B(N2027), .Y(N2070) );
  NOR2X1 gate587 ( .A(N2028), .B(N2029), .Y(N2073) );
  NOR2X1 gate588 ( .A(N2030), .B(N1176), .Y(N2076) );
  NOR2X1 gate589 ( .A(N2001), .B(N2033), .Y(N2080) );
  NOR2X1 gate590 ( .A(N2033), .B(N1224), .Y(N2081) );
  NOR2X1 gate591 ( .A(N1897), .B(N2033), .Y(N2082) );
  NOR2X1 gate592 ( .A(N2037), .B(N552), .Y(N2085) );
  NOR2X1 gate593 ( .A(N2040), .B(N600), .Y(N2089) );
  NOR2X1 gate594 ( .A(N2043), .B(N648), .Y(N2093) );
  NOR2X1 gate595 ( .A(N2046), .B(N696), .Y(N2097) );
  NOR2X1 gate596 ( .A(N2049), .B(N744), .Y(N2101) );
  NOR2X1 gate597 ( .A(N2052), .B(N792), .Y(N2105) );
  NOR2X1 gate598 ( .A(N2055), .B(N840), .Y(N2109) );
  NOR2X1 gate599 ( .A(N2058), .B(N888), .Y(N2113) );
  NOR2X1 gate600 ( .A(N2061), .B(N936), .Y(N2117) );
  NOR2X1 gate601 ( .A(N2064), .B(N984), .Y(N2121) );
  NOR2X1 gate602 ( .A(N2067), .B(N1032), .Y(N2125) );
  NOR2X1 gate603 ( .A(N2070), .B(N1080), .Y(N2129) );
  NOR2X1 gate604 ( .A(N2073), .B(N1128), .Y(N2133) );
  NOR2X1 gate605 ( .A(N2030), .B(N2076), .Y(N2137) );
  NOR2X1 gate606 ( .A(N2076), .B(N1176), .Y(N2138) );
  NOR2X1 gate607 ( .A(N1941), .B(N2076), .Y(N2139) );
  NOR2X1 gate608 ( .A(N2080), .B(N2081), .Y(N2142) );
  NOR2X1 gate609 ( .A(N1272), .B(N2082), .Y(N2145) );
  NOR2X1 gate610 ( .A(N2037), .B(N2085), .Y(N2149) );
  NOR2X1 gate611 ( .A(N2085), .B(N552), .Y(N2150) );
  NOR2X1 gate612 ( .A(N1947), .B(N2085), .Y(N2151) );
  NOR2X1 gate613 ( .A(N2040), .B(N2089), .Y(N2154) );
  NOR2X1 gate614 ( .A(N2089), .B(N600), .Y(N2155) );
  NOR2X1 gate615 ( .A(N1951), .B(N2089), .Y(N2156) );
  NOR2X1 gate616 ( .A(N2043), .B(N2093), .Y(N2159) );
  NOR2X1 gate617 ( .A(N2093), .B(N648), .Y(N2160) );
  NOR2X1 gate618 ( .A(N1955), .B(N2093), .Y(N2161) );
  NOR2X1 gate619 ( .A(N2046), .B(N2097), .Y(N2164) );
  NOR2X1 gate620 ( .A(N2097), .B(N696), .Y(N2165) );
  NOR2X1 gate621 ( .A(N1959), .B(N2097), .Y(N2166) );
  NOR2X1 gate622 ( .A(N2049), .B(N2101), .Y(N2169) );
  NOR2X1 gate623 ( .A(N2101), .B(N744), .Y(N2170) );
  NOR2X1 gate624 ( .A(N1963), .B(N2101), .Y(N2171) );
  NOR2X1 gate625 ( .A(N2052), .B(N2105), .Y(N2174) );
  NOR2X1 gate626 ( .A(N2105), .B(N792), .Y(N2175) );
  NOR2X1 gate627 ( .A(N1967), .B(N2105), .Y(N2176) );
  NOR2X1 gate628 ( .A(N2055), .B(N2109), .Y(N2179) );
  NOR2X1 gate629 ( .A(N2109), .B(N840), .Y(N2180) );
  NOR2X1 gate630 ( .A(N1971), .B(N2109), .Y(N2181) );
  NOR2X1 gate631 ( .A(N2058), .B(N2113), .Y(N2184) );
  NOR2X1 gate632 ( .A(N2113), .B(N888), .Y(N2185) );
  NOR2X1 gate633 ( .A(N1975), .B(N2113), .Y(N2186) );
  NOR2X1 gate634 ( .A(N2061), .B(N2117), .Y(N2189) );
  NOR2X1 gate635 ( .A(N2117), .B(N936), .Y(N2190) );
  NOR2X1 gate636 ( .A(N1979), .B(N2117), .Y(N2191) );
  NOR2X1 gate637 ( .A(N2064), .B(N2121), .Y(N2194) );
  NOR2X1 gate638 ( .A(N2121), .B(N984), .Y(N2195) );
  NOR2X1 gate639 ( .A(N1983), .B(N2121), .Y(N2196) );
  NOR2X1 gate640 ( .A(N2067), .B(N2125), .Y(N2199) );
  NOR2X1 gate641 ( .A(N2125), .B(N1032), .Y(N2200) );
  NOR2X1 gate642 ( .A(N1987), .B(N2125), .Y(N2201) );
  NOR2X1 gate643 ( .A(N2070), .B(N2129), .Y(N2204) );
  NOR2X1 gate644 ( .A(N2129), .B(N1080), .Y(N2205) );
  NOR2X1 gate645 ( .A(N1991), .B(N2129), .Y(N2206) );
  NOR2X1 gate646 ( .A(N2073), .B(N2133), .Y(N2209) );
  NOR2X1 gate647 ( .A(N2133), .B(N1128), .Y(N2210) );
  NOR2X1 gate648 ( .A(N1995), .B(N2133), .Y(N2211) );
  NOR2X1 gate649 ( .A(N2137), .B(N2138), .Y(N2214) );
  NOR2X1 gate650 ( .A(N2142), .B(N2139), .Y(N2217) );
  NOR2X1 gate651 ( .A(N1272), .B(N2145), .Y(N2221) );
  NOR2X1 gate652 ( .A(N2145), .B(N2082), .Y(N2222) );
  NOR2X1 gate653 ( .A(N2149), .B(N2150), .Y(N2223) );
  NOR2X1 gate654 ( .A(N2154), .B(N2155), .Y(N2224) );
  NOR2X1 gate655 ( .A(N2159), .B(N2160), .Y(N2227) );
  NOR2X1 gate656 ( .A(N2164), .B(N2165), .Y(N2230) );
  NOR2X1 gate657 ( .A(N2169), .B(N2170), .Y(N2233) );
  NOR2X1 gate658 ( .A(N2174), .B(N2175), .Y(N2236) );
  NOR2X1 gate659 ( .A(N2179), .B(N2180), .Y(N2239) );
  NOR2X1 gate660 ( .A(N2184), .B(N2185), .Y(N2242) );
  NOR2X1 gate661 ( .A(N2189), .B(N2190), .Y(N2245) );
  NOR2X1 gate662 ( .A(N2194), .B(N2195), .Y(N2248) );
  NOR2X1 gate663 ( .A(N2199), .B(N2200), .Y(N2251) );
  NOR2X1 gate664 ( .A(N2204), .B(N2205), .Y(N2254) );
  NOR2X1 gate665 ( .A(N2209), .B(N2210), .Y(N2257) );
  NOR2X1 gate666 ( .A(N2214), .B(N2211), .Y(N2260) );
  NOR2X1 gate667 ( .A(N2142), .B(N2217), .Y(N2264) );
  NOR2X1 gate668 ( .A(N2217), .B(N2139), .Y(N2265) );
  NOR2X1 gate669 ( .A(N2221), .B(N2222), .Y(N2266) );
  NOR2X1 gate670 ( .A(N2224), .B(N2151), .Y(N2269) );
  NOR2X1 gate671 ( .A(N2227), .B(N2156), .Y(N2273) );
  NOR2X1 gate672 ( .A(N2230), .B(N2161), .Y(N2277) );
  NOR2X1 gate673 ( .A(N2233), .B(N2166), .Y(N2281) );
  NOR2X1 gate674 ( .A(N2236), .B(N2171), .Y(N2285) );
  NOR2X1 gate675 ( .A(N2239), .B(N2176), .Y(N2289) );
  NOR2X1 gate676 ( .A(N2242), .B(N2181), .Y(N2293) );
  NOR2X1 gate677 ( .A(N2245), .B(N2186), .Y(N2297) );
  NOR2X1 gate678 ( .A(N2248), .B(N2191), .Y(N2301) );
  NOR2X1 gate679 ( .A(N2251), .B(N2196), .Y(N2305) );
  NOR2X1 gate680 ( .A(N2254), .B(N2201), .Y(N2309) );
  NOR2X1 gate681 ( .A(N2257), .B(N2206), .Y(N2313) );
  NOR2X1 gate682 ( .A(N2214), .B(N2260), .Y(N2317) );
  NOR2X1 gate683 ( .A(N2260), .B(N2211), .Y(N2318) );
  NOR2X1 gate684 ( .A(N2264), .B(N2265), .Y(N2319) );
  NOR2X1 gate685 ( .A(N2266), .B(N1227), .Y(N2322) );
  NOR2X1 gate686 ( .A(N2224), .B(N2269), .Y(N2326) );
  NOR2X1 gate687 ( .A(N2269), .B(N2151), .Y(N2327) );
  NOR2X1 gate688 ( .A(N2227), .B(N2273), .Y(N2328) );
  NOR2X1 gate689 ( .A(N2273), .B(N2156), .Y(N2329) );
  NOR2X1 gate690 ( .A(N2230), .B(N2277), .Y(N2330) );
  NOR2X1 gate691 ( .A(N2277), .B(N2161), .Y(N2331) );
  NOR2X1 gate692 ( .A(N2233), .B(N2281), .Y(N2332) );
  NOR2X1 gate693 ( .A(N2281), .B(N2166), .Y(N2333) );
  NOR2X1 gate694 ( .A(N2236), .B(N2285), .Y(N2334) );
  NOR2X1 gate695 ( .A(N2285), .B(N2171), .Y(N2335) );
  NOR2X1 gate696 ( .A(N2239), .B(N2289), .Y(N2336) );
  NOR2X1 gate697 ( .A(N2289), .B(N2176), .Y(N2337) );
  NOR2X1 gate698 ( .A(N2242), .B(N2293), .Y(N2338) );
  NOR2X1 gate699 ( .A(N2293), .B(N2181), .Y(N2339) );
  NOR2X1 gate700 ( .A(N2245), .B(N2297), .Y(N2340) );
  NOR2X1 gate701 ( .A(N2297), .B(N2186), .Y(N2341) );
  NOR2X1 gate702 ( .A(N2248), .B(N2301), .Y(N2342) );
  NOR2X1 gate703 ( .A(N2301), .B(N2191), .Y(N2343) );
  NOR2X1 gate704 ( .A(N2251), .B(N2305), .Y(N2344) );
  NOR2X1 gate705 ( .A(N2305), .B(N2196), .Y(N2345) );
  NOR2X1 gate706 ( .A(N2254), .B(N2309), .Y(N2346) );
  NOR2X1 gate707 ( .A(N2309), .B(N2201), .Y(N2347) );
  NOR2X1 gate708 ( .A(N2257), .B(N2313), .Y(N2348) );
  NOR2X1 gate709 ( .A(N2313), .B(N2206), .Y(N2349) );
  NOR2X1 gate710 ( .A(N2317), .B(N2318), .Y(N2350) );
  NOR2X1 gate711 ( .A(N2319), .B(N1179), .Y(N2353) );
  NOR2X1 gate712 ( .A(N2266), .B(N2322), .Y(N2357) );
  NOR2X1 gate713 ( .A(N2322), .B(N1227), .Y(N2358) );
  NOR2X1 gate714 ( .A(N2145), .B(N2322), .Y(N2359) );
  NOR2X1 gate715 ( .A(N2326), .B(N2327), .Y(N2362) );
  NOR2X1 gate716 ( .A(N2328), .B(N2329), .Y(N2365) );
  NOR2X1 gate717 ( .A(N2330), .B(N2331), .Y(N2368) );
  NOR2X1 gate718 ( .A(N2332), .B(N2333), .Y(N2371) );
  NOR2X1 gate719 ( .A(N2334), .B(N2335), .Y(N2374) );
  NOR2X1 gate720 ( .A(N2336), .B(N2337), .Y(N2377) );
  NOR2X1 gate721 ( .A(N2338), .B(N2339), .Y(N2380) );
  NOR2X1 gate722 ( .A(N2340), .B(N2341), .Y(N2383) );
  NOR2X1 gate723 ( .A(N2342), .B(N2343), .Y(N2386) );
  NOR2X1 gate724 ( .A(N2344), .B(N2345), .Y(N2389) );
  NOR2X1 gate725 ( .A(N2346), .B(N2347), .Y(N2392) );
  NOR2X1 gate726 ( .A(N2348), .B(N2349), .Y(N2395) );
  NOR2X1 gate727 ( .A(N2350), .B(N1131), .Y(N2398) );
  NOR2X1 gate728 ( .A(N2319), .B(N2353), .Y(N2402) );
  NOR2X1 gate729 ( .A(N2353), .B(N1179), .Y(N2403) );
  NOR2X1 gate730 ( .A(N2217), .B(N2353), .Y(N2404) );
  NOR2X1 gate731 ( .A(N2357), .B(N2358), .Y(N2407) );
  NOR2X1 gate732 ( .A(N1275), .B(N2359), .Y(N2410) );
  NOR2X1 gate733 ( .A(N2362), .B(N555), .Y(N2414) );
  NOR2X1 gate734 ( .A(N2365), .B(N603), .Y(N2418) );
  NOR2X1 gate735 ( .A(N2368), .B(N651), .Y(N2422) );
  NOR2X1 gate736 ( .A(N2371), .B(N699), .Y(N2426) );
  NOR2X1 gate737 ( .A(N2374), .B(N747), .Y(N2430) );
  NOR2X1 gate738 ( .A(N2377), .B(N795), .Y(N2434) );
  NOR2X1 gate739 ( .A(N2380), .B(N843), .Y(N2438) );
  NOR2X1 gate740 ( .A(N2383), .B(N891), .Y(N2442) );
  NOR2X1 gate741 ( .A(N2386), .B(N939), .Y(N2446) );
  NOR2X1 gate742 ( .A(N2389), .B(N987), .Y(N2450) );
  NOR2X1 gate743 ( .A(N2392), .B(N1035), .Y(N2454) );
  NOR2X1 gate744 ( .A(N2395), .B(N1083), .Y(N2458) );
  NOR2X1 gate745 ( .A(N2350), .B(N2398), .Y(N2462) );
  NOR2X1 gate746 ( .A(N2398), .B(N1131), .Y(N2463) );
  NOR2X1 gate747 ( .A(N2260), .B(N2398), .Y(N2464) );
  NOR2X1 gate748 ( .A(N2402), .B(N2403), .Y(N2467) );
  NOR2X1 gate749 ( .A(N2407), .B(N2404), .Y(N2470) );
  NOR2X1 gate750 ( .A(N1275), .B(N2410), .Y(N2474) );
  NOR2X1 gate751 ( .A(N2410), .B(N2359), .Y(N2475) );
  NOR2X1 gate752 ( .A(N2362), .B(N2414), .Y(N2476) );
  NOR2X1 gate753 ( .A(N2414), .B(N555), .Y(N2477) );
  NOR2X1 gate754 ( .A(N2269), .B(N2414), .Y(N2478) );
  NOR2X1 gate755 ( .A(N2365), .B(N2418), .Y(N2481) );
  NOR2X1 gate756 ( .A(N2418), .B(N603), .Y(N2482) );
  NOR2X1 gate757 ( .A(N2273), .B(N2418), .Y(N2483) );
  NOR2X1 gate758 ( .A(N2368), .B(N2422), .Y(N2486) );
  NOR2X1 gate759 ( .A(N2422), .B(N651), .Y(N2487) );
  NOR2X1 gate760 ( .A(N2277), .B(N2422), .Y(N2488) );
  NOR2X1 gate761 ( .A(N2371), .B(N2426), .Y(N2491) );
  NOR2X1 gate762 ( .A(N2426), .B(N699), .Y(N2492) );
  NOR2X1 gate763 ( .A(N2281), .B(N2426), .Y(N2493) );
  NOR2X1 gate764 ( .A(N2374), .B(N2430), .Y(N2496) );
  NOR2X1 gate765 ( .A(N2430), .B(N747), .Y(N2497) );
  NOR2X1 gate766 ( .A(N2285), .B(N2430), .Y(N2498) );
  NOR2X1 gate767 ( .A(N2377), .B(N2434), .Y(N2501) );
  NOR2X1 gate768 ( .A(N2434), .B(N795), .Y(N2502) );
  NOR2X1 gate769 ( .A(N2289), .B(N2434), .Y(N2503) );
  NOR2X1 gate770 ( .A(N2380), .B(N2438), .Y(N2506) );
  NOR2X1 gate771 ( .A(N2438), .B(N843), .Y(N2507) );
  NOR2X1 gate772 ( .A(N2293), .B(N2438), .Y(N2508) );
  NOR2X1 gate773 ( .A(N2383), .B(N2442), .Y(N2511) );
  NOR2X1 gate774 ( .A(N2442), .B(N891), .Y(N2512) );
  NOR2X1 gate775 ( .A(N2297), .B(N2442), .Y(N2513) );
  NOR2X1 gate776 ( .A(N2386), .B(N2446), .Y(N2516) );
  NOR2X1 gate777 ( .A(N2446), .B(N939), .Y(N2517) );
  NOR2X1 gate778 ( .A(N2301), .B(N2446), .Y(N2518) );
  NOR2X1 gate779 ( .A(N2389), .B(N2450), .Y(N2521) );
  NOR2X1 gate780 ( .A(N2450), .B(N987), .Y(N2522) );
  NOR2X1 gate781 ( .A(N2305), .B(N2450), .Y(N2523) );
  NOR2X1 gate782 ( .A(N2392), .B(N2454), .Y(N2526) );
  NOR2X1 gate783 ( .A(N2454), .B(N1035), .Y(N2527) );
  NOR2X1 gate784 ( .A(N2309), .B(N2454), .Y(N2528) );
  NOR2X1 gate785 ( .A(N2395), .B(N2458), .Y(N2531) );
  NOR2X1 gate786 ( .A(N2458), .B(N1083), .Y(N2532) );
  NOR2X1 gate787 ( .A(N2313), .B(N2458), .Y(N2533) );
  NOR2X1 gate788 ( .A(N2462), .B(N2463), .Y(N2536) );
  NOR2X1 gate789 ( .A(N2467), .B(N2464), .Y(N2539) );
  NOR2X1 gate790 ( .A(N2407), .B(N2470), .Y(N2543) );
  NOR2X1 gate791 ( .A(N2470), .B(N2404), .Y(N2544) );
  NOR2X1 gate792 ( .A(N2474), .B(N2475), .Y(N2545) );
  NOR2X1 gate793 ( .A(N2476), .B(N2477), .Y(N2548) );
  NOR2X1 gate794 ( .A(N2481), .B(N2482), .Y(N2549) );
  NOR2X1 gate795 ( .A(N2486), .B(N2487), .Y(N2552) );
  NOR2X1 gate796 ( .A(N2491), .B(N2492), .Y(N2555) );
  NOR2X1 gate797 ( .A(N2496), .B(N2497), .Y(N2558) );
  NOR2X1 gate798 ( .A(N2501), .B(N2502), .Y(N2561) );
  NOR2X1 gate799 ( .A(N2506), .B(N2507), .Y(N2564) );
  NOR2X1 gate800 ( .A(N2511), .B(N2512), .Y(N2567) );
  NOR2X1 gate801 ( .A(N2516), .B(N2517), .Y(N2570) );
  NOR2X1 gate802 ( .A(N2521), .B(N2522), .Y(N2573) );
  NOR2X1 gate803 ( .A(N2526), .B(N2527), .Y(N2576) );
  NOR2X1 gate804 ( .A(N2531), .B(N2532), .Y(N2579) );
  NOR2X1 gate805 ( .A(N2536), .B(N2533), .Y(N2582) );
  NOR2X1 gate806 ( .A(N2467), .B(N2539), .Y(N2586) );
  NOR2X1 gate807 ( .A(N2539), .B(N2464), .Y(N2587) );
  NOR2X1 gate808 ( .A(N2543), .B(N2544), .Y(N2588) );
  NOR2X1 gate809 ( .A(N2545), .B(N1230), .Y(N2591) );
  NOR2X1 gate810 ( .A(N2549), .B(N2478), .Y(N2595) );
  NOR2X1 gate811 ( .A(N2552), .B(N2483), .Y(N2599) );
  NOR2X1 gate812 ( .A(N2555), .B(N2488), .Y(N2603) );
  NOR2X1 gate813 ( .A(N2558), .B(N2493), .Y(N2607) );
  NOR2X1 gate814 ( .A(N2561), .B(N2498), .Y(N2611) );
  NOR2X1 gate815 ( .A(N2564), .B(N2503), .Y(N2615) );
  NOR2X1 gate816 ( .A(N2567), .B(N2508), .Y(N2619) );
  NOR2X1 gate817 ( .A(N2570), .B(N2513), .Y(N2623) );
  NOR2X1 gate818 ( .A(N2573), .B(N2518), .Y(N2627) );
  NOR2X1 gate819 ( .A(N2576), .B(N2523), .Y(N2631) );
  NOR2X1 gate820 ( .A(N2579), .B(N2528), .Y(N2635) );
  NOR2X1 gate821 ( .A(N2536), .B(N2582), .Y(N2639) );
  NOR2X1 gate822 ( .A(N2582), .B(N2533), .Y(N2640) );
  NOR2X1 gate823 ( .A(N2586), .B(N2587), .Y(N2641) );
  NOR2X1 gate824 ( .A(N2588), .B(N1182), .Y(N2644) );
  NOR2X1 gate825 ( .A(N2545), .B(N2591), .Y(N2648) );
  NOR2X1 gate826 ( .A(N2591), .B(N1230), .Y(N2649) );
  NOR2X1 gate827 ( .A(N2410), .B(N2591), .Y(N2650) );
  NOR2X1 gate828 ( .A(N2549), .B(N2595), .Y(N2653) );
  NOR2X1 gate829 ( .A(N2595), .B(N2478), .Y(N2654) );
  NOR2X1 gate830 ( .A(N2552), .B(N2599), .Y(N2655) );
  NOR2X1 gate831 ( .A(N2599), .B(N2483), .Y(N2656) );
  NOR2X1 gate832 ( .A(N2555), .B(N2603), .Y(N2657) );
  NOR2X1 gate833 ( .A(N2603), .B(N2488), .Y(N2658) );
  NOR2X1 gate834 ( .A(N2558), .B(N2607), .Y(N2659) );
  NOR2X1 gate835 ( .A(N2607), .B(N2493), .Y(N2660) );
  NOR2X1 gate836 ( .A(N2561), .B(N2611), .Y(N2661) );
  NOR2X1 gate837 ( .A(N2611), .B(N2498), .Y(N2662) );
  NOR2X1 gate838 ( .A(N2564), .B(N2615), .Y(N2663) );
  NOR2X1 gate839 ( .A(N2615), .B(N2503), .Y(N2664) );
  NOR2X1 gate840 ( .A(N2567), .B(N2619), .Y(N2665) );
  NOR2X1 gate841 ( .A(N2619), .B(N2508), .Y(N2666) );
  NOR2X1 gate842 ( .A(N2570), .B(N2623), .Y(N2667) );
  NOR2X1 gate843 ( .A(N2623), .B(N2513), .Y(N2668) );
  NOR2X1 gate844 ( .A(N2573), .B(N2627), .Y(N2669) );
  NOR2X1 gate845 ( .A(N2627), .B(N2518), .Y(N2670) );
  NOR2X1 gate846 ( .A(N2576), .B(N2631), .Y(N2671) );
  NOR2X1 gate847 ( .A(N2631), .B(N2523), .Y(N2672) );
  NOR2X1 gate848 ( .A(N2579), .B(N2635), .Y(N2673) );
  NOR2X1 gate849 ( .A(N2635), .B(N2528), .Y(N2674) );
  NOR2X1 gate850 ( .A(N2639), .B(N2640), .Y(N2675) );
  NOR2X1 gate851 ( .A(N2641), .B(N1134), .Y(N2678) );
  NOR2X1 gate852 ( .A(N2588), .B(N2644), .Y(N2682) );
  NOR2X1 gate853 ( .A(N2644), .B(N1182), .Y(N2683) );
  NOR2X1 gate854 ( .A(N2470), .B(N2644), .Y(N2684) );
  NOR2X1 gate855 ( .A(N2648), .B(N2649), .Y(N2687) );
  NOR2X1 gate856 ( .A(N1278), .B(N2650), .Y(N2690) );
  NOR2X1 gate857 ( .A(N2653), .B(N2654), .Y(N2694) );
  NOR2X1 gate858 ( .A(N2655), .B(N2656), .Y(N2697) );
  NOR2X1 gate859 ( .A(N2657), .B(N2658), .Y(N2700) );
  NOR2X1 gate860 ( .A(N2659), .B(N2660), .Y(N2703) );
  NOR2X1 gate861 ( .A(N2661), .B(N2662), .Y(N2706) );
  NOR2X1 gate862 ( .A(N2663), .B(N2664), .Y(N2709) );
  NOR2X1 gate863 ( .A(N2665), .B(N2666), .Y(N2712) );
  NOR2X1 gate864 ( .A(N2667), .B(N2668), .Y(N2715) );
  NOR2X1 gate865 ( .A(N2669), .B(N2670), .Y(N2718) );
  NOR2X1 gate866 ( .A(N2671), .B(N2672), .Y(N2721) );
  NOR2X1 gate867 ( .A(N2673), .B(N2674), .Y(N2724) );
  NOR2X1 gate868 ( .A(N2675), .B(N1086), .Y(N2727) );
  NOR2X1 gate869 ( .A(N2641), .B(N2678), .Y(N2731) );
  NOR2X1 gate870 ( .A(N2678), .B(N1134), .Y(N2732) );
  NOR2X1 gate871 ( .A(N2539), .B(N2678), .Y(N2733) );
  NOR2X1 gate872 ( .A(N2682), .B(N2683), .Y(N2736) );
  NOR2X1 gate873 ( .A(N2687), .B(N2684), .Y(N2739) );
  NOR2X1 gate874 ( .A(N1278), .B(N2690), .Y(N2743) );
  NOR2X1 gate875 ( .A(N2690), .B(N2650), .Y(N2744) );
  NOR2X1 gate876 ( .A(N2694), .B(N558), .Y(N2745) );
  NOR2X1 gate877 ( .A(N2697), .B(N606), .Y(N2749) );
  NOR2X1 gate878 ( .A(N2700), .B(N654), .Y(N2753) );
  NOR2X1 gate879 ( .A(N2703), .B(N702), .Y(N2757) );
  NOR2X1 gate880 ( .A(N2706), .B(N750), .Y(N2761) );
  NOR2X1 gate881 ( .A(N2709), .B(N798), .Y(N2765) );
  NOR2X1 gate882 ( .A(N2712), .B(N846), .Y(N2769) );
  NOR2X1 gate883 ( .A(N2715), .B(N894), .Y(N2773) );
  NOR2X1 gate884 ( .A(N2718), .B(N942), .Y(N2777) );
  NOR2X1 gate885 ( .A(N2721), .B(N990), .Y(N2781) );
  NOR2X1 gate886 ( .A(N2724), .B(N1038), .Y(N2785) );
  NOR2X1 gate887 ( .A(N2675), .B(N2727), .Y(N2789) );
  NOR2X1 gate888 ( .A(N2727), .B(N1086), .Y(N2790) );
  NOR2X1 gate889 ( .A(N2582), .B(N2727), .Y(N2791) );
  NOR2X1 gate890 ( .A(N2731), .B(N2732), .Y(N2794) );
  NOR2X1 gate891 ( .A(N2736), .B(N2733), .Y(N2797) );
  NOR2X1 gate892 ( .A(N2687), .B(N2739), .Y(N2801) );
  NOR2X1 gate893 ( .A(N2739), .B(N2684), .Y(N2802) );
  NOR2X1 gate894 ( .A(N2743), .B(N2744), .Y(N2803) );
  NOR2X1 gate895 ( .A(N2694), .B(N2745), .Y(N2806) );
  NOR2X1 gate896 ( .A(N2745), .B(N558), .Y(N2807) );
  NOR2X1 gate897 ( .A(N2595), .B(N2745), .Y(N2808) );
  NOR2X1 gate898 ( .A(N2697), .B(N2749), .Y(N2811) );
  NOR2X1 gate899 ( .A(N2749), .B(N606), .Y(N2812) );
  NOR2X1 gate900 ( .A(N2599), .B(N2749), .Y(N2813) );
  NOR2X1 gate901 ( .A(N2700), .B(N2753), .Y(N2816) );
  NOR2X1 gate902 ( .A(N2753), .B(N654), .Y(N2817) );
  NOR2X1 gate903 ( .A(N2603), .B(N2753), .Y(N2818) );
  NOR2X1 gate904 ( .A(N2703), .B(N2757), .Y(N2821) );
  NOR2X1 gate905 ( .A(N2757), .B(N702), .Y(N2822) );
  NOR2X1 gate906 ( .A(N2607), .B(N2757), .Y(N2823) );
  NOR2X1 gate907 ( .A(N2706), .B(N2761), .Y(N2826) );
  NOR2X1 gate908 ( .A(N2761), .B(N750), .Y(N2827) );
  NOR2X1 gate909 ( .A(N2611), .B(N2761), .Y(N2828) );
  NOR2X1 gate910 ( .A(N2709), .B(N2765), .Y(N2831) );
  NOR2X1 gate911 ( .A(N2765), .B(N798), .Y(N2832) );
  NOR2X1 gate912 ( .A(N2615), .B(N2765), .Y(N2833) );
  NOR2X1 gate913 ( .A(N2712), .B(N2769), .Y(N2836) );
  NOR2X1 gate914 ( .A(N2769), .B(N846), .Y(N2837) );
  NOR2X1 gate915 ( .A(N2619), .B(N2769), .Y(N2838) );
  NOR2X1 gate916 ( .A(N2715), .B(N2773), .Y(N2841) );
  NOR2X1 gate917 ( .A(N2773), .B(N894), .Y(N2842) );
  NOR2X1 gate918 ( .A(N2623), .B(N2773), .Y(N2843) );
  NOR2X1 gate919 ( .A(N2718), .B(N2777), .Y(N2846) );
  NOR2X1 gate920 ( .A(N2777), .B(N942), .Y(N2847) );
  NOR2X1 gate921 ( .A(N2627), .B(N2777), .Y(N2848) );
  NOR2X1 gate922 ( .A(N2721), .B(N2781), .Y(N2851) );
  NOR2X1 gate923 ( .A(N2781), .B(N990), .Y(N2852) );
  NOR2X1 gate924 ( .A(N2631), .B(N2781), .Y(N2853) );
  NOR2X1 gate925 ( .A(N2724), .B(N2785), .Y(N2856) );
  NOR2X1 gate926 ( .A(N2785), .B(N1038), .Y(N2857) );
  NOR2X1 gate927 ( .A(N2635), .B(N2785), .Y(N2858) );
  NOR2X1 gate928 ( .A(N2789), .B(N2790), .Y(N2861) );
  NOR2X1 gate929 ( .A(N2794), .B(N2791), .Y(N2864) );
  NOR2X1 gate930 ( .A(N2736), .B(N2797), .Y(N2868) );
  NOR2X1 gate931 ( .A(N2797), .B(N2733), .Y(N2869) );
  NOR2X1 gate932 ( .A(N2801), .B(N2802), .Y(N2870) );
  NOR2X1 gate933 ( .A(N2803), .B(N1233), .Y(N2873) );
  NOR2X1 gate934 ( .A(N2806), .B(N2807), .Y(N2877) );
  NOR2X1 gate935 ( .A(N2811), .B(N2812), .Y(N2878) );
  NOR2X1 gate936 ( .A(N2816), .B(N2817), .Y(N2881) );
  NOR2X1 gate937 ( .A(N2821), .B(N2822), .Y(N2884) );
  NOR2X1 gate938 ( .A(N2826), .B(N2827), .Y(N2887) );
  NOR2X1 gate939 ( .A(N2831), .B(N2832), .Y(N2890) );
  NOR2X1 gate940 ( .A(N2836), .B(N2837), .Y(N2893) );
  NOR2X1 gate941 ( .A(N2841), .B(N2842), .Y(N2896) );
  NOR2X1 gate942 ( .A(N2846), .B(N2847), .Y(N2899) );
  NOR2X1 gate943 ( .A(N2851), .B(N2852), .Y(N2902) );
  NOR2X1 gate944 ( .A(N2856), .B(N2857), .Y(N2905) );
  NOR2X1 gate945 ( .A(N2861), .B(N2858), .Y(N2908) );
  NOR2X1 gate946 ( .A(N2794), .B(N2864), .Y(N2912) );
  NOR2X1 gate947 ( .A(N2864), .B(N2791), .Y(N2913) );
  NOR2X1 gate948 ( .A(N2868), .B(N2869), .Y(N2914) );
  NOR2X1 gate949 ( .A(N2870), .B(N1185), .Y(N2917) );
  NOR2X1 gate950 ( .A(N2803), .B(N2873), .Y(N2921) );
  NOR2X1 gate951 ( .A(N2873), .B(N1233), .Y(N2922) );
  NOR2X1 gate952 ( .A(N2690), .B(N2873), .Y(N2923) );
  NOR2X1 gate953 ( .A(N2878), .B(N2808), .Y(N2926) );
  NOR2X1 gate954 ( .A(N2881), .B(N2813), .Y(N2930) );
  NOR2X1 gate955 ( .A(N2884), .B(N2818), .Y(N2934) );
  NOR2X1 gate956 ( .A(N2887), .B(N2823), .Y(N2938) );
  NOR2X1 gate957 ( .A(N2890), .B(N2828), .Y(N2942) );
  NOR2X1 gate958 ( .A(N2893), .B(N2833), .Y(N2946) );
  NOR2X1 gate959 ( .A(N2896), .B(N2838), .Y(N2950) );
  NOR2X1 gate960 ( .A(N2899), .B(N2843), .Y(N2954) );
  NOR2X1 gate961 ( .A(N2902), .B(N2848), .Y(N2958) );
  NOR2X1 gate962 ( .A(N2905), .B(N2853), .Y(N2962) );
  NOR2X1 gate963 ( .A(N2861), .B(N2908), .Y(N2966) );
  NOR2X1 gate964 ( .A(N2908), .B(N2858), .Y(N2967) );
  NOR2X1 gate965 ( .A(N2912), .B(N2913), .Y(N2968) );
  NOR2X1 gate966 ( .A(N2914), .B(N1137), .Y(N2971) );
  NOR2X1 gate967 ( .A(N2870), .B(N2917), .Y(N2975) );
  NOR2X1 gate968 ( .A(N2917), .B(N1185), .Y(N2976) );
  NOR2X1 gate969 ( .A(N2739), .B(N2917), .Y(N2977) );
  NOR2X1 gate970 ( .A(N2921), .B(N2922), .Y(N2980) );
  NOR2X1 gate971 ( .A(N1281), .B(N2923), .Y(N2983) );
  NOR2X1 gate972 ( .A(N2878), .B(N2926), .Y(N2987) );
  NOR2X1 gate973 ( .A(N2926), .B(N2808), .Y(N2988) );
  NOR2X1 gate974 ( .A(N2881), .B(N2930), .Y(N2989) );
  NOR2X1 gate975 ( .A(N2930), .B(N2813), .Y(N2990) );
  NOR2X1 gate976 ( .A(N2884), .B(N2934), .Y(N2991) );
  NOR2X1 gate977 ( .A(N2934), .B(N2818), .Y(N2992) );
  NOR2X1 gate978 ( .A(N2887), .B(N2938), .Y(N2993) );
  NOR2X1 gate979 ( .A(N2938), .B(N2823), .Y(N2994) );
  NOR2X1 gate980 ( .A(N2890), .B(N2942), .Y(N2995) );
  NOR2X1 gate981 ( .A(N2942), .B(N2828), .Y(N2996) );
  NOR2X1 gate982 ( .A(N2893), .B(N2946), .Y(N2997) );
  NOR2X1 gate983 ( .A(N2946), .B(N2833), .Y(N2998) );
  NOR2X1 gate984 ( .A(N2896), .B(N2950), .Y(N2999) );
  NOR2X1 gate985 ( .A(N2950), .B(N2838), .Y(N3000) );
  NOR2X1 gate986 ( .A(N2899), .B(N2954), .Y(N3001) );
  NOR2X1 gate987 ( .A(N2954), .B(N2843), .Y(N3002) );
  NOR2X1 gate988 ( .A(N2902), .B(N2958), .Y(N3003) );
  NOR2X1 gate989 ( .A(N2958), .B(N2848), .Y(N3004) );
  NOR2X1 gate990 ( .A(N2905), .B(N2962), .Y(N3005) );
  NOR2X1 gate991 ( .A(N2962), .B(N2853), .Y(N3006) );
  NOR2X1 gate992 ( .A(N2966), .B(N2967), .Y(N3007) );
  NOR2X1 gate993 ( .A(N2968), .B(N1089), .Y(N3010) );
  NOR2X1 gate994 ( .A(N2914), .B(N2971), .Y(N3014) );
  NOR2X1 gate995 ( .A(N2971), .B(N1137), .Y(N3015) );
  NOR2X1 gate996 ( .A(N2797), .B(N2971), .Y(N3016) );
  NOR2X1 gate997 ( .A(N2975), .B(N2976), .Y(N3019) );
  NOR2X1 gate998 ( .A(N2980), .B(N2977), .Y(N3022) );
  NOR2X1 gate999 ( .A(N1281), .B(N2983), .Y(N3026) );
  NOR2X1 gate1000 ( .A(N2983), .B(N2923), .Y(N3027) );
  NOR2X1 gate1001 ( .A(N2987), .B(N2988), .Y(N3028) );
  NOR2X1 gate1002 ( .A(N2989), .B(N2990), .Y(N3031) );
  NOR2X1 gate1003 ( .A(N2991), .B(N2992), .Y(N3034) );
  NOR2X1 gate1004 ( .A(N2993), .B(N2994), .Y(N3037) );
  NOR2X1 gate1005 ( .A(N2995), .B(N2996), .Y(N3040) );
  NOR2X1 gate1006 ( .A(N2997), .B(N2998), .Y(N3043) );
  NOR2X1 gate1007 ( .A(N2999), .B(N3000), .Y(N3046) );
  NOR2X1 gate1008 ( .A(N3001), .B(N3002), .Y(N3049) );
  NOR2X1 gate1009 ( .A(N3003), .B(N3004), .Y(N3052) );
  NOR2X1 gate1010 ( .A(N3005), .B(N3006), .Y(N3055) );
  NOR2X1 gate1011 ( .A(N3007), .B(N1041), .Y(N3058) );
  NOR2X1 gate1012 ( .A(N2968), .B(N3010), .Y(N3062) );
  NOR2X1 gate1013 ( .A(N3010), .B(N1089), .Y(N3063) );
  NOR2X1 gate1014 ( .A(N2864), .B(N3010), .Y(N3064) );
  NOR2X1 gate1015 ( .A(N3014), .B(N3015), .Y(N3067) );
  NOR2X1 gate1016 ( .A(N3019), .B(N3016), .Y(N3070) );
  NOR2X1 gate1017 ( .A(N2980), .B(N3022), .Y(N3074) );
  NOR2X1 gate1018 ( .A(N3022), .B(N2977), .Y(N3075) );
  NOR2X1 gate1019 ( .A(N3026), .B(N3027), .Y(N3076) );
  NOR2X1 gate1020 ( .A(N3028), .B(N561), .Y(N3079) );
  NOR2X1 gate1021 ( .A(N3031), .B(N609), .Y(N3083) );
  NOR2X1 gate1022 ( .A(N3034), .B(N657), .Y(N3087) );
  NOR2X1 gate1023 ( .A(N3037), .B(N705), .Y(N3091) );
  NOR2X1 gate1024 ( .A(N3040), .B(N753), .Y(N3095) );
  NOR2X1 gate1025 ( .A(N3043), .B(N801), .Y(N3099) );
  NOR2X1 gate1026 ( .A(N3046), .B(N849), .Y(N3103) );
  NOR2X1 gate1027 ( .A(N3049), .B(N897), .Y(N3107) );
  NOR2X1 gate1028 ( .A(N3052), .B(N945), .Y(N3111) );
  NOR2X1 gate1029 ( .A(N3055), .B(N993), .Y(N3115) );
  NOR2X1 gate1030 ( .A(N3007), .B(N3058), .Y(N3119) );
  NOR2X1 gate1031 ( .A(N3058), .B(N1041), .Y(N3120) );
  NOR2X1 gate1032 ( .A(N2908), .B(N3058), .Y(N3121) );
  NOR2X1 gate1033 ( .A(N3062), .B(N3063), .Y(N3124) );
  NOR2X1 gate1034 ( .A(N3067), .B(N3064), .Y(N3127) );
  NOR2X1 gate1035 ( .A(N3019), .B(N3070), .Y(N3131) );
  NOR2X1 gate1036 ( .A(N3070), .B(N3016), .Y(N3132) );
  NOR2X1 gate1037 ( .A(N3074), .B(N3075), .Y(N3133) );
  NOR2X1 gate1038 ( .A(N3076), .B(N1236), .Y(N3136) );
  NOR2X1 gate1039 ( .A(N3028), .B(N3079), .Y(N3140) );
  NOR2X1 gate1040 ( .A(N3079), .B(N561), .Y(N3141) );
  NOR2X1 gate1041 ( .A(N2926), .B(N3079), .Y(N3142) );
  NOR2X1 gate1042 ( .A(N3031), .B(N3083), .Y(N3145) );
  NOR2X1 gate1043 ( .A(N3083), .B(N609), .Y(N3146) );
  NOR2X1 gate1044 ( .A(N2930), .B(N3083), .Y(N3147) );
  NOR2X1 gate1045 ( .A(N3034), .B(N3087), .Y(N3150) );
  NOR2X1 gate1046 ( .A(N3087), .B(N657), .Y(N3151) );
  NOR2X1 gate1047 ( .A(N2934), .B(N3087), .Y(N3152) );
  NOR2X1 gate1048 ( .A(N3037), .B(N3091), .Y(N3155) );
  NOR2X1 gate1049 ( .A(N3091), .B(N705), .Y(N3156) );
  NOR2X1 gate1050 ( .A(N2938), .B(N3091), .Y(N3157) );
  NOR2X1 gate1051 ( .A(N3040), .B(N3095), .Y(N3160) );
  NOR2X1 gate1052 ( .A(N3095), .B(N753), .Y(N3161) );
  NOR2X1 gate1053 ( .A(N2942), .B(N3095), .Y(N3162) );
  NOR2X1 gate1054 ( .A(N3043), .B(N3099), .Y(N3165) );
  NOR2X1 gate1055 ( .A(N3099), .B(N801), .Y(N3166) );
  NOR2X1 gate1056 ( .A(N2946), .B(N3099), .Y(N3167) );
  NOR2X1 gate1057 ( .A(N3046), .B(N3103), .Y(N3170) );
  NOR2X1 gate1058 ( .A(N3103), .B(N849), .Y(N3171) );
  NOR2X1 gate1059 ( .A(N2950), .B(N3103), .Y(N3172) );
  NOR2X1 gate1060 ( .A(N3049), .B(N3107), .Y(N3175) );
  NOR2X1 gate1061 ( .A(N3107), .B(N897), .Y(N3176) );
  NOR2X1 gate1062 ( .A(N2954), .B(N3107), .Y(N3177) );
  NOR2X1 gate1063 ( .A(N3052), .B(N3111), .Y(N3180) );
  NOR2X1 gate1064 ( .A(N3111), .B(N945), .Y(N3181) );
  NOR2X1 gate1065 ( .A(N2958), .B(N3111), .Y(N3182) );
  NOR2X1 gate1066 ( .A(N3055), .B(N3115), .Y(N3185) );
  NOR2X1 gate1067 ( .A(N3115), .B(N993), .Y(N3186) );
  NOR2X1 gate1068 ( .A(N2962), .B(N3115), .Y(N3187) );
  NOR2X1 gate1069 ( .A(N3119), .B(N3120), .Y(N3190) );
  NOR2X1 gate1070 ( .A(N3124), .B(N3121), .Y(N3193) );
  NOR2X1 gate1071 ( .A(N3067), .B(N3127), .Y(N3197) );
  NOR2X1 gate1072 ( .A(N3127), .B(N3064), .Y(N3198) );
  NOR2X1 gate1073 ( .A(N3131), .B(N3132), .Y(N3199) );
  NOR2X1 gate1074 ( .A(N3133), .B(N1188), .Y(N3202) );
  NOR2X1 gate1075 ( .A(N3076), .B(N3136), .Y(N3206) );
  NOR2X1 gate1076 ( .A(N3136), .B(N1236), .Y(N3207) );
  NOR2X1 gate1077 ( .A(N2983), .B(N3136), .Y(N3208) );
  NOR2X1 gate1078 ( .A(N3140), .B(N3141), .Y(N3211) );
  NOR2X1 gate1079 ( .A(N3145), .B(N3146), .Y(N3212) );
  NOR2X1 gate1080 ( .A(N3150), .B(N3151), .Y(N3215) );
  NOR2X1 gate1081 ( .A(N3155), .B(N3156), .Y(N3218) );
  NOR2X1 gate1082 ( .A(N3160), .B(N3161), .Y(N3221) );
  NOR2X1 gate1083 ( .A(N3165), .B(N3166), .Y(N3224) );
  NOR2X1 gate1084 ( .A(N3170), .B(N3171), .Y(N3227) );
  NOR2X1 gate1085 ( .A(N3175), .B(N3176), .Y(N3230) );
  NOR2X1 gate1086 ( .A(N3180), .B(N3181), .Y(N3233) );
  NOR2X1 gate1087 ( .A(N3185), .B(N3186), .Y(N3236) );
  NOR2X1 gate1088 ( .A(N3190), .B(N3187), .Y(N3239) );
  NOR2X1 gate1089 ( .A(N3124), .B(N3193), .Y(N3243) );
  NOR2X1 gate1090 ( .A(N3193), .B(N3121), .Y(N3244) );
  NOR2X1 gate1091 ( .A(N3197), .B(N3198), .Y(N3245) );
  NOR2X1 gate1092 ( .A(N3199), .B(N1140), .Y(N3248) );
  NOR2X1 gate1093 ( .A(N3133), .B(N3202), .Y(N3252) );
  NOR2X1 gate1094 ( .A(N3202), .B(N1188), .Y(N3253) );
  NOR2X1 gate1095 ( .A(N3022), .B(N3202), .Y(N3254) );
  NOR2X1 gate1096 ( .A(N3206), .B(N3207), .Y(N3257) );
  NOR2X1 gate1097 ( .A(N1284), .B(N3208), .Y(N3260) );
  NOR2X1 gate1098 ( .A(N3212), .B(N3142), .Y(N3264) );
  NOR2X1 gate1099 ( .A(N3215), .B(N3147), .Y(N3268) );
  NOR2X1 gate1100 ( .A(N3218), .B(N3152), .Y(N3272) );
  NOR2X1 gate1101 ( .A(N3221), .B(N3157), .Y(N3276) );
  NOR2X1 gate1102 ( .A(N3224), .B(N3162), .Y(N3280) );
  NOR2X1 gate1103 ( .A(N3227), .B(N3167), .Y(N3284) );
  NOR2X1 gate1104 ( .A(N3230), .B(N3172), .Y(N3288) );
  NOR2X1 gate1105 ( .A(N3233), .B(N3177), .Y(N3292) );
  NOR2X1 gate1106 ( .A(N3236), .B(N3182), .Y(N3296) );
  NOR2X1 gate1107 ( .A(N3190), .B(N3239), .Y(N3300) );
  NOR2X1 gate1108 ( .A(N3239), .B(N3187), .Y(N3301) );
  NOR2X1 gate1109 ( .A(N3243), .B(N3244), .Y(N3302) );
  NOR2X1 gate1110 ( .A(N3245), .B(N1092), .Y(N3305) );
  NOR2X1 gate1111 ( .A(N3199), .B(N3248), .Y(N3309) );
  NOR2X1 gate1112 ( .A(N3248), .B(N1140), .Y(N3310) );
  NOR2X1 gate1113 ( .A(N3070), .B(N3248), .Y(N3311) );
  NOR2X1 gate1114 ( .A(N3252), .B(N3253), .Y(N3314) );
  NOR2X1 gate1115 ( .A(N3257), .B(N3254), .Y(N3317) );
  NOR2X1 gate1116 ( .A(N1284), .B(N3260), .Y(N3321) );
  NOR2X1 gate1117 ( .A(N3260), .B(N3208), .Y(N3322) );
  NOR2X1 gate1118 ( .A(N3212), .B(N3264), .Y(N3323) );
  NOR2X1 gate1119 ( .A(N3264), .B(N3142), .Y(N3324) );
  NOR2X1 gate1120 ( .A(N3215), .B(N3268), .Y(N3325) );
  NOR2X1 gate1121 ( .A(N3268), .B(N3147), .Y(N3326) );
  NOR2X1 gate1122 ( .A(N3218), .B(N3272), .Y(N3327) );
  NOR2X1 gate1123 ( .A(N3272), .B(N3152), .Y(N3328) );
  NOR2X1 gate1124 ( .A(N3221), .B(N3276), .Y(N3329) );
  NOR2X1 gate1125 ( .A(N3276), .B(N3157), .Y(N3330) );
  NOR2X1 gate1126 ( .A(N3224), .B(N3280), .Y(N3331) );
  NOR2X1 gate1127 ( .A(N3280), .B(N3162), .Y(N3332) );
  NOR2X1 gate1128 ( .A(N3227), .B(N3284), .Y(N3333) );
  NOR2X1 gate1129 ( .A(N3284), .B(N3167), .Y(N3334) );
  NOR2X1 gate1130 ( .A(N3230), .B(N3288), .Y(N3335) );
  NOR2X1 gate1131 ( .A(N3288), .B(N3172), .Y(N3336) );
  NOR2X1 gate1132 ( .A(N3233), .B(N3292), .Y(N3337) );
  NOR2X1 gate1133 ( .A(N3292), .B(N3177), .Y(N3338) );
  NOR2X1 gate1134 ( .A(N3236), .B(N3296), .Y(N3339) );
  NOR2X1 gate1135 ( .A(N3296), .B(N3182), .Y(N3340) );
  NOR2X1 gate1136 ( .A(N3300), .B(N3301), .Y(N3341) );
  NOR2X1 gate1137 ( .A(N3302), .B(N1044), .Y(N3344) );
  NOR2X1 gate1138 ( .A(N3245), .B(N3305), .Y(N3348) );
  NOR2X1 gate1139 ( .A(N3305), .B(N1092), .Y(N3349) );
  NOR2X1 gate1140 ( .A(N3127), .B(N3305), .Y(N3350) );
  NOR2X1 gate1141 ( .A(N3309), .B(N3310), .Y(N3353) );
  NOR2X1 gate1142 ( .A(N3314), .B(N3311), .Y(N3356) );
  NOR2X1 gate1143 ( .A(N3257), .B(N3317), .Y(N3360) );
  NOR2X1 gate1144 ( .A(N3317), .B(N3254), .Y(N3361) );
  NOR2X1 gate1145 ( .A(N3321), .B(N3322), .Y(N3362) );
  NOR2X1 gate1146 ( .A(N3323), .B(N3324), .Y(N3365) );
  NOR2X1 gate1147 ( .A(N3325), .B(N3326), .Y(N3368) );
  NOR2X1 gate1148 ( .A(N3327), .B(N3328), .Y(N3371) );
  NOR2X1 gate1149 ( .A(N3329), .B(N3330), .Y(N3374) );
  NOR2X1 gate1150 ( .A(N3331), .B(N3332), .Y(N3377) );
  NOR2X1 gate1151 ( .A(N3333), .B(N3334), .Y(N3380) );
  NOR2X1 gate1152 ( .A(N3335), .B(N3336), .Y(N3383) );
  NOR2X1 gate1153 ( .A(N3337), .B(N3338), .Y(N3386) );
  NOR2X1 gate1154 ( .A(N3339), .B(N3340), .Y(N3389) );
  NOR2X1 gate1155 ( .A(N3341), .B(N996), .Y(N3392) );
  NOR2X1 gate1156 ( .A(N3302), .B(N3344), .Y(N3396) );
  NOR2X1 gate1157 ( .A(N3344), .B(N1044), .Y(N3397) );
  NOR2X1 gate1158 ( .A(N3193), .B(N3344), .Y(N3398) );
  NOR2X1 gate1159 ( .A(N3348), .B(N3349), .Y(N3401) );
  NOR2X1 gate1160 ( .A(N3353), .B(N3350), .Y(N3404) );
  NOR2X1 gate1161 ( .A(N3314), .B(N3356), .Y(N3408) );
  NOR2X1 gate1162 ( .A(N3356), .B(N3311), .Y(N3409) );
  NOR2X1 gate1163 ( .A(N3360), .B(N3361), .Y(N3410) );
  NOR2X1 gate1164 ( .A(N3362), .B(N1239), .Y(N3413) );
  NOR2X1 gate1165 ( .A(N3365), .B(N564), .Y(N3417) );
  NOR2X1 gate1166 ( .A(N3368), .B(N612), .Y(N3421) );
  NOR2X1 gate1167 ( .A(N3371), .B(N660), .Y(N3425) );
  NOR2X1 gate1168 ( .A(N3374), .B(N708), .Y(N3429) );
  NOR2X1 gate1169 ( .A(N3377), .B(N756), .Y(N3433) );
  NOR2X1 gate1170 ( .A(N3380), .B(N804), .Y(N3437) );
  NOR2X1 gate1171 ( .A(N3383), .B(N852), .Y(N3441) );
  NOR2X1 gate1172 ( .A(N3386), .B(N900), .Y(N3445) );
  NOR2X1 gate1173 ( .A(N3389), .B(N948), .Y(N3449) );
  NOR2X1 gate1174 ( .A(N3341), .B(N3392), .Y(N3453) );
  NOR2X1 gate1175 ( .A(N3392), .B(N996), .Y(N3454) );
  NOR2X1 gate1176 ( .A(N3239), .B(N3392), .Y(N3455) );
  NOR2X1 gate1177 ( .A(N3396), .B(N3397), .Y(N3458) );
  NOR2X1 gate1178 ( .A(N3401), .B(N3398), .Y(N3461) );
  NOR2X1 gate1179 ( .A(N3353), .B(N3404), .Y(N3465) );
  NOR2X1 gate1180 ( .A(N3404), .B(N3350), .Y(N3466) );
  NOR2X1 gate1181 ( .A(N3408), .B(N3409), .Y(N3467) );
  NOR2X1 gate1182 ( .A(N3410), .B(N1191), .Y(N3470) );
  NOR2X1 gate1183 ( .A(N3362), .B(N3413), .Y(N3474) );
  NOR2X1 gate1184 ( .A(N3413), .B(N1239), .Y(N3475) );
  NOR2X1 gate1185 ( .A(N3260), .B(N3413), .Y(N3476) );
  NOR2X1 gate1186 ( .A(N3365), .B(N3417), .Y(N3479) );
  NOR2X1 gate1187 ( .A(N3417), .B(N564), .Y(N3480) );
  NOR2X1 gate1188 ( .A(N3264), .B(N3417), .Y(N3481) );
  NOR2X1 gate1189 ( .A(N3368), .B(N3421), .Y(N3484) );
  NOR2X1 gate1190 ( .A(N3421), .B(N612), .Y(N3485) );
  NOR2X1 gate1191 ( .A(N3268), .B(N3421), .Y(N3486) );
  NOR2X1 gate1192 ( .A(N3371), .B(N3425), .Y(N3489) );
  NOR2X1 gate1193 ( .A(N3425), .B(N660), .Y(N3490) );
  NOR2X1 gate1194 ( .A(N3272), .B(N3425), .Y(N3491) );
  NOR2X1 gate1195 ( .A(N3374), .B(N3429), .Y(N3494) );
  NOR2X1 gate1196 ( .A(N3429), .B(N708), .Y(N3495) );
  NOR2X1 gate1197 ( .A(N3276), .B(N3429), .Y(N3496) );
  NOR2X1 gate1198 ( .A(N3377), .B(N3433), .Y(N3499) );
  NOR2X1 gate1199 ( .A(N3433), .B(N756), .Y(N3500) );
  NOR2X1 gate1200 ( .A(N3280), .B(N3433), .Y(N3501) );
  NOR2X1 gate1201 ( .A(N3380), .B(N3437), .Y(N3504) );
  NOR2X1 gate1202 ( .A(N3437), .B(N804), .Y(N3505) );
  NOR2X1 gate1203 ( .A(N3284), .B(N3437), .Y(N3506) );
  NOR2X1 gate1204 ( .A(N3383), .B(N3441), .Y(N3509) );
  NOR2X1 gate1205 ( .A(N3441), .B(N852), .Y(N3510) );
  NOR2X1 gate1206 ( .A(N3288), .B(N3441), .Y(N3511) );
  NOR2X1 gate1207 ( .A(N3386), .B(N3445), .Y(N3514) );
  NOR2X1 gate1208 ( .A(N3445), .B(N900), .Y(N3515) );
  NOR2X1 gate1209 ( .A(N3292), .B(N3445), .Y(N3516) );
  NOR2X1 gate1210 ( .A(N3389), .B(N3449), .Y(N3519) );
  NOR2X1 gate1211 ( .A(N3449), .B(N948), .Y(N3520) );
  NOR2X1 gate1212 ( .A(N3296), .B(N3449), .Y(N3521) );
  NOR2X1 gate1213 ( .A(N3453), .B(N3454), .Y(N3524) );
  NOR2X1 gate1214 ( .A(N3458), .B(N3455), .Y(N3527) );
  NOR2X1 gate1215 ( .A(N3401), .B(N3461), .Y(N3531) );
  NOR2X1 gate1216 ( .A(N3461), .B(N3398), .Y(N3532) );
  NOR2X1 gate1217 ( .A(N3465), .B(N3466), .Y(N3533) );
  NOR2X1 gate1218 ( .A(N3467), .B(N1143), .Y(N3536) );
  NOR2X1 gate1219 ( .A(N3410), .B(N3470), .Y(N3540) );
  NOR2X1 gate1220 ( .A(N3470), .B(N1191), .Y(N3541) );
  NOR2X1 gate1221 ( .A(N3317), .B(N3470), .Y(N3542) );
  NOR2X1 gate1222 ( .A(N3474), .B(N3475), .Y(N3545) );
  NOR2X1 gate1223 ( .A(N1287), .B(N3476), .Y(N3548) );
  NOR2X1 gate1224 ( .A(N3479), .B(N3480), .Y(N3552) );
  NOR2X1 gate1225 ( .A(N3484), .B(N3485), .Y(N3553) );
  NOR2X1 gate1226 ( .A(N3489), .B(N3490), .Y(N3556) );
  NOR2X1 gate1227 ( .A(N3494), .B(N3495), .Y(N3559) );
  NOR2X1 gate1228 ( .A(N3499), .B(N3500), .Y(N3562) );
  NOR2X1 gate1229 ( .A(N3504), .B(N3505), .Y(N3565) );
  NOR2X1 gate1230 ( .A(N3509), .B(N3510), .Y(N3568) );
  NOR2X1 gate1231 ( .A(N3514), .B(N3515), .Y(N3571) );
  NOR2X1 gate1232 ( .A(N3519), .B(N3520), .Y(N3574) );
  NOR2X1 gate1233 ( .A(N3524), .B(N3521), .Y(N3577) );
  NOR2X1 gate1234 ( .A(N3458), .B(N3527), .Y(N3581) );
  NOR2X1 gate1235 ( .A(N3527), .B(N3455), .Y(N3582) );
  NOR2X1 gate1236 ( .A(N3531), .B(N3532), .Y(N3583) );
  NOR2X1 gate1237 ( .A(N3533), .B(N1095), .Y(N3586) );
  NOR2X1 gate1238 ( .A(N3467), .B(N3536), .Y(N3590) );
  NOR2X1 gate1239 ( .A(N3536), .B(N1143), .Y(N3591) );
  NOR2X1 gate1240 ( .A(N3356), .B(N3536), .Y(N3592) );
  NOR2X1 gate1241 ( .A(N3540), .B(N3541), .Y(N3595) );
  NOR2X1 gate1242 ( .A(N3545), .B(N3542), .Y(N3598) );
  NOR2X1 gate1243 ( .A(N1287), .B(N3548), .Y(N3602) );
  NOR2X1 gate1244 ( .A(N3548), .B(N3476), .Y(N3603) );
  NOR2X1 gate1245 ( .A(N3553), .B(N3481), .Y(N3604) );
  NOR2X1 gate1246 ( .A(N3556), .B(N3486), .Y(N3608) );
  NOR2X1 gate1247 ( .A(N3559), .B(N3491), .Y(N3612) );
  NOR2X1 gate1248 ( .A(N3562), .B(N3496), .Y(N3616) );
  NOR2X1 gate1249 ( .A(N3565), .B(N3501), .Y(N3620) );
  NOR2X1 gate1250 ( .A(N3568), .B(N3506), .Y(N3624) );
  NOR2X1 gate1251 ( .A(N3571), .B(N3511), .Y(N3628) );
  NOR2X1 gate1252 ( .A(N3574), .B(N3516), .Y(N3632) );
  NOR2X1 gate1253 ( .A(N3524), .B(N3577), .Y(N3636) );
  NOR2X1 gate1254 ( .A(N3577), .B(N3521), .Y(N3637) );
  NOR2X1 gate1255 ( .A(N3581), .B(N3582), .Y(N3638) );
  NOR2X1 gate1256 ( .A(N3583), .B(N1047), .Y(N3641) );
  NOR2X1 gate1257 ( .A(N3533), .B(N3586), .Y(N3645) );
  NOR2X1 gate1258 ( .A(N3586), .B(N1095), .Y(N3646) );
  NOR2X1 gate1259 ( .A(N3404), .B(N3586), .Y(N3647) );
  NOR2X1 gate1260 ( .A(N3590), .B(N3591), .Y(N3650) );
  NOR2X1 gate1261 ( .A(N3595), .B(N3592), .Y(N3653) );
  NOR2X1 gate1262 ( .A(N3545), .B(N3598), .Y(N3657) );
  NOR2X1 gate1263 ( .A(N3598), .B(N3542), .Y(N3658) );
  NOR2X1 gate1264 ( .A(N3602), .B(N3603), .Y(N3659) );
  NOR2X1 gate1265 ( .A(N3553), .B(N3604), .Y(N3662) );
  NOR2X1 gate1266 ( .A(N3604), .B(N3481), .Y(N3663) );
  NOR2X1 gate1267 ( .A(N3556), .B(N3608), .Y(N3664) );
  NOR2X1 gate1268 ( .A(N3608), .B(N3486), .Y(N3665) );
  NOR2X1 gate1269 ( .A(N3559), .B(N3612), .Y(N3666) );
  NOR2X1 gate1270 ( .A(N3612), .B(N3491), .Y(N3667) );
  NOR2X1 gate1271 ( .A(N3562), .B(N3616), .Y(N3668) );
  NOR2X1 gate1272 ( .A(N3616), .B(N3496), .Y(N3669) );
  NOR2X1 gate1273 ( .A(N3565), .B(N3620), .Y(N3670) );
  NOR2X1 gate1274 ( .A(N3620), .B(N3501), .Y(N3671) );
  NOR2X1 gate1275 ( .A(N3568), .B(N3624), .Y(N3672) );
  NOR2X1 gate1276 ( .A(N3624), .B(N3506), .Y(N3673) );
  NOR2X1 gate1277 ( .A(N3571), .B(N3628), .Y(N3674) );
  NOR2X1 gate1278 ( .A(N3628), .B(N3511), .Y(N3675) );
  NOR2X1 gate1279 ( .A(N3574), .B(N3632), .Y(N3676) );
  NOR2X1 gate1280 ( .A(N3632), .B(N3516), .Y(N3677) );
  NOR2X1 gate1281 ( .A(N3636), .B(N3637), .Y(N3678) );
  NOR2X1 gate1282 ( .A(N3638), .B(N999), .Y(N3681) );
  NOR2X1 gate1283 ( .A(N3583), .B(N3641), .Y(N3685) );
  NOR2X1 gate1284 ( .A(N3641), .B(N1047), .Y(N3686) );
  NOR2X1 gate1285 ( .A(N3461), .B(N3641), .Y(N3687) );
  NOR2X1 gate1286 ( .A(N3645), .B(N3646), .Y(N3690) );
  NOR2X1 gate1287 ( .A(N3650), .B(N3647), .Y(N3693) );
  NOR2X1 gate1288 ( .A(N3595), .B(N3653), .Y(N3697) );
  NOR2X1 gate1289 ( .A(N3653), .B(N3592), .Y(N3698) );
  NOR2X1 gate1290 ( .A(N3657), .B(N3658), .Y(N3699) );
  NOR2X1 gate1291 ( .A(N3659), .B(N1242), .Y(N3702) );
  NOR2X1 gate1292 ( .A(N3662), .B(N3663), .Y(N3706) );
  NOR2X1 gate1293 ( .A(N3664), .B(N3665), .Y(N3709) );
  NOR2X1 gate1294 ( .A(N3666), .B(N3667), .Y(N3712) );
  NOR2X1 gate1295 ( .A(N3668), .B(N3669), .Y(N3715) );
  NOR2X1 gate1296 ( .A(N3670), .B(N3671), .Y(N3718) );
  NOR2X1 gate1297 ( .A(N3672), .B(N3673), .Y(N3721) );
  NOR2X1 gate1298 ( .A(N3674), .B(N3675), .Y(N3724) );
  NOR2X1 gate1299 ( .A(N3676), .B(N3677), .Y(N3727) );
  NOR2X1 gate1300 ( .A(N3678), .B(N951), .Y(N3730) );
  NOR2X1 gate1301 ( .A(N3638), .B(N3681), .Y(N3734) );
  NOR2X1 gate1302 ( .A(N3681), .B(N999), .Y(N3735) );
  NOR2X1 gate1303 ( .A(N3527), .B(N3681), .Y(N3736) );
  NOR2X1 gate1304 ( .A(N3685), .B(N3686), .Y(N3739) );
  NOR2X1 gate1305 ( .A(N3690), .B(N3687), .Y(N3742) );
  NOR2X1 gate1306 ( .A(N3650), .B(N3693), .Y(N3746) );
  NOR2X1 gate1307 ( .A(N3693), .B(N3647), .Y(N3747) );
  NOR2X1 gate1308 ( .A(N3697), .B(N3698), .Y(N3748) );
  NOR2X1 gate1309 ( .A(N3699), .B(N1194), .Y(N3751) );
  NOR2X1 gate1310 ( .A(N3659), .B(N3702), .Y(N3755) );
  NOR2X1 gate1311 ( .A(N3702), .B(N1242), .Y(N3756) );
  NOR2X1 gate1312 ( .A(N3548), .B(N3702), .Y(N3757) );
  NOR2X1 gate1313 ( .A(N3706), .B(N567), .Y(N3760) );
  NOR2X1 gate1314 ( .A(N3709), .B(N615), .Y(N3764) );
  NOR2X1 gate1315 ( .A(N3712), .B(N663), .Y(N3768) );
  NOR2X1 gate1316 ( .A(N3715), .B(N711), .Y(N3772) );
  NOR2X1 gate1317 ( .A(N3718), .B(N759), .Y(N3776) );
  NOR2X1 gate1318 ( .A(N3721), .B(N807), .Y(N3780) );
  NOR2X1 gate1319 ( .A(N3724), .B(N855), .Y(N3784) );
  NOR2X1 gate1320 ( .A(N3727), .B(N903), .Y(N3788) );
  NOR2X1 gate1321 ( .A(N3678), .B(N3730), .Y(N3792) );
  NOR2X1 gate1322 ( .A(N3730), .B(N951), .Y(N3793) );
  NOR2X1 gate1323 ( .A(N3577), .B(N3730), .Y(N3794) );
  NOR2X1 gate1324 ( .A(N3734), .B(N3735), .Y(N3797) );
  NOR2X1 gate1325 ( .A(N3739), .B(N3736), .Y(N3800) );
  NOR2X1 gate1326 ( .A(N3690), .B(N3742), .Y(N3804) );
  NOR2X1 gate1327 ( .A(N3742), .B(N3687), .Y(N3805) );
  NOR2X1 gate1328 ( .A(N3746), .B(N3747), .Y(N3806) );
  NOR2X1 gate1329 ( .A(N3748), .B(N1146), .Y(N3809) );
  NOR2X1 gate1330 ( .A(N3699), .B(N3751), .Y(N3813) );
  NOR2X1 gate1331 ( .A(N3751), .B(N1194), .Y(N3814) );
  NOR2X1 gate1332 ( .A(N3598), .B(N3751), .Y(N3815) );
  NOR2X1 gate1333 ( .A(N3755), .B(N3756), .Y(N3818) );
  NOR2X1 gate1334 ( .A(N1290), .B(N3757), .Y(N3821) );
  NOR2X1 gate1335 ( .A(N3706), .B(N3760), .Y(N3825) );
  NOR2X1 gate1336 ( .A(N3760), .B(N567), .Y(N3826) );
  NOR2X1 gate1337 ( .A(N3604), .B(N3760), .Y(N3827) );
  NOR2X1 gate1338 ( .A(N3709), .B(N3764), .Y(N3830) );
  NOR2X1 gate1339 ( .A(N3764), .B(N615), .Y(N3831) );
  NOR2X1 gate1340 ( .A(N3608), .B(N3764), .Y(N3832) );
  NOR2X1 gate1341 ( .A(N3712), .B(N3768), .Y(N3835) );
  NOR2X1 gate1342 ( .A(N3768), .B(N663), .Y(N3836) );
  NOR2X1 gate1343 ( .A(N3612), .B(N3768), .Y(N3837) );
  NOR2X1 gate1344 ( .A(N3715), .B(N3772), .Y(N3840) );
  NOR2X1 gate1345 ( .A(N3772), .B(N711), .Y(N3841) );
  NOR2X1 gate1346 ( .A(N3616), .B(N3772), .Y(N3842) );
  NOR2X1 gate1347 ( .A(N3718), .B(N3776), .Y(N3845) );
  NOR2X1 gate1348 ( .A(N3776), .B(N759), .Y(N3846) );
  NOR2X1 gate1349 ( .A(N3620), .B(N3776), .Y(N3847) );
  NOR2X1 gate1350 ( .A(N3721), .B(N3780), .Y(N3850) );
  NOR2X1 gate1351 ( .A(N3780), .B(N807), .Y(N3851) );
  NOR2X1 gate1352 ( .A(N3624), .B(N3780), .Y(N3852) );
  NOR2X1 gate1353 ( .A(N3724), .B(N3784), .Y(N3855) );
  NOR2X1 gate1354 ( .A(N3784), .B(N855), .Y(N3856) );
  NOR2X1 gate1355 ( .A(N3628), .B(N3784), .Y(N3857) );
  NOR2X1 gate1356 ( .A(N3727), .B(N3788), .Y(N3860) );
  NOR2X1 gate1357 ( .A(N3788), .B(N903), .Y(N3861) );
  NOR2X1 gate1358 ( .A(N3632), .B(N3788), .Y(N3862) );
  NOR2X1 gate1359 ( .A(N3792), .B(N3793), .Y(N3865) );
  NOR2X1 gate1360 ( .A(N3797), .B(N3794), .Y(N3868) );
  NOR2X1 gate1361 ( .A(N3739), .B(N3800), .Y(N3872) );
  NOR2X1 gate1362 ( .A(N3800), .B(N3736), .Y(N3873) );
  NOR2X1 gate1363 ( .A(N3804), .B(N3805), .Y(N3874) );
  NOR2X1 gate1364 ( .A(N3806), .B(N1098), .Y(N3877) );
  NOR2X1 gate1365 ( .A(N3748), .B(N3809), .Y(N3881) );
  NOR2X1 gate1366 ( .A(N3809), .B(N1146), .Y(N3882) );
  NOR2X1 gate1367 ( .A(N3653), .B(N3809), .Y(N3883) );
  NOR2X1 gate1368 ( .A(N3813), .B(N3814), .Y(N3886) );
  NOR2X1 gate1369 ( .A(N3818), .B(N3815), .Y(N3889) );
  NOR2X1 gate1370 ( .A(N1290), .B(N3821), .Y(N3893) );
  NOR2X1 gate1371 ( .A(N3821), .B(N3757), .Y(N3894) );
  NOR2X1 gate1372 ( .A(N3825), .B(N3826), .Y(N3895) );
  NOR2X1 gate1373 ( .A(N3830), .B(N3831), .Y(N3896) );
  NOR2X1 gate1374 ( .A(N3835), .B(N3836), .Y(N3899) );
  NOR2X1 gate1375 ( .A(N3840), .B(N3841), .Y(N3902) );
  NOR2X1 gate1376 ( .A(N3845), .B(N3846), .Y(N3905) );
  NOR2X1 gate1377 ( .A(N3850), .B(N3851), .Y(N3908) );
  NOR2X1 gate1378 ( .A(N3855), .B(N3856), .Y(N3911) );
  NOR2X1 gate1379 ( .A(N3860), .B(N3861), .Y(N3914) );
  NOR2X1 gate1380 ( .A(N3865), .B(N3862), .Y(N3917) );
  NOR2X1 gate1381 ( .A(N3797), .B(N3868), .Y(N3921) );
  NOR2X1 gate1382 ( .A(N3868), .B(N3794), .Y(N3922) );
  NOR2X1 gate1383 ( .A(N3872), .B(N3873), .Y(N3923) );
  NOR2X1 gate1384 ( .A(N3874), .B(N1050), .Y(N3926) );
  NOR2X1 gate1385 ( .A(N3806), .B(N3877), .Y(N3930) );
  NOR2X1 gate1386 ( .A(N3877), .B(N1098), .Y(N3931) );
  NOR2X1 gate1387 ( .A(N3693), .B(N3877), .Y(N3932) );
  NOR2X1 gate1388 ( .A(N3881), .B(N3882), .Y(N3935) );
  NOR2X1 gate1389 ( .A(N3886), .B(N3883), .Y(N3938) );
  NOR2X1 gate1390 ( .A(N3818), .B(N3889), .Y(N3942) );
  NOR2X1 gate1391 ( .A(N3889), .B(N3815), .Y(N3943) );
  NOR2X1 gate1392 ( .A(N3893), .B(N3894), .Y(N3944) );
  NOR2X1 gate1393 ( .A(N3896), .B(N3827), .Y(N3947) );
  NOR2X1 gate1394 ( .A(N3899), .B(N3832), .Y(N3951) );
  NOR2X1 gate1395 ( .A(N3902), .B(N3837), .Y(N3955) );
  NOR2X1 gate1396 ( .A(N3905), .B(N3842), .Y(N3959) );
  NOR2X1 gate1397 ( .A(N3908), .B(N3847), .Y(N3963) );
  NOR2X1 gate1398 ( .A(N3911), .B(N3852), .Y(N3967) );
  NOR2X1 gate1399 ( .A(N3914), .B(N3857), .Y(N3971) );
  NOR2X1 gate1400 ( .A(N3865), .B(N3917), .Y(N3975) );
  NOR2X1 gate1401 ( .A(N3917), .B(N3862), .Y(N3976) );
  NOR2X1 gate1402 ( .A(N3921), .B(N3922), .Y(N3977) );
  NOR2X1 gate1403 ( .A(N3923), .B(N1002), .Y(N3980) );
  NOR2X1 gate1404 ( .A(N3874), .B(N3926), .Y(N3984) );
  NOR2X1 gate1405 ( .A(N3926), .B(N1050), .Y(N3985) );
  NOR2X1 gate1406 ( .A(N3742), .B(N3926), .Y(N3986) );
  NOR2X1 gate1407 ( .A(N3930), .B(N3931), .Y(N3989) );
  NOR2X1 gate1408 ( .A(N3935), .B(N3932), .Y(N3992) );
  NOR2X1 gate1409 ( .A(N3886), .B(N3938), .Y(N3996) );
  NOR2X1 gate1410 ( .A(N3938), .B(N3883), .Y(N3997) );
  NOR2X1 gate1411 ( .A(N3942), .B(N3943), .Y(N3998) );
  NOR2X1 gate1412 ( .A(N3944), .B(N1245), .Y(N4001) );
  NOR2X1 gate1413 ( .A(N3896), .B(N3947), .Y(N4005) );
  NOR2X1 gate1414 ( .A(N3947), .B(N3827), .Y(N4006) );
  NOR2X1 gate1415 ( .A(N3899), .B(N3951), .Y(N4007) );
  NOR2X1 gate1416 ( .A(N3951), .B(N3832), .Y(N4008) );
  NOR2X1 gate1417 ( .A(N3902), .B(N3955), .Y(N4009) );
  NOR2X1 gate1418 ( .A(N3955), .B(N3837), .Y(N4010) );
  NOR2X1 gate1419 ( .A(N3905), .B(N3959), .Y(N4011) );
  NOR2X1 gate1420 ( .A(N3959), .B(N3842), .Y(N4012) );
  NOR2X1 gate1421 ( .A(N3908), .B(N3963), .Y(N4013) );
  NOR2X1 gate1422 ( .A(N3963), .B(N3847), .Y(N4014) );
  NOR2X1 gate1423 ( .A(N3911), .B(N3967), .Y(N4015) );
  NOR2X1 gate1424 ( .A(N3967), .B(N3852), .Y(N4016) );
  NOR2X1 gate1425 ( .A(N3914), .B(N3971), .Y(N4017) );
  NOR2X1 gate1426 ( .A(N3971), .B(N3857), .Y(N4018) );
  NOR2X1 gate1427 ( .A(N3975), .B(N3976), .Y(N4019) );
  NOR2X1 gate1428 ( .A(N3977), .B(N954), .Y(N4022) );
  NOR2X1 gate1429 ( .A(N3923), .B(N3980), .Y(N4026) );
  NOR2X1 gate1430 ( .A(N3980), .B(N1002), .Y(N4027) );
  NOR2X1 gate1431 ( .A(N3800), .B(N3980), .Y(N4028) );
  NOR2X1 gate1432 ( .A(N3984), .B(N3985), .Y(N4031) );
  NOR2X1 gate1433 ( .A(N3989), .B(N3986), .Y(N4034) );
  NOR2X1 gate1434 ( .A(N3935), .B(N3992), .Y(N4038) );
  NOR2X1 gate1435 ( .A(N3992), .B(N3932), .Y(N4039) );
  NOR2X1 gate1436 ( .A(N3996), .B(N3997), .Y(N4040) );
  NOR2X1 gate1437 ( .A(N3998), .B(N1197), .Y(N4043) );
  NOR2X1 gate1438 ( .A(N3944), .B(N4001), .Y(N4047) );
  NOR2X1 gate1439 ( .A(N4001), .B(N1245), .Y(N4048) );
  NOR2X1 gate1440 ( .A(N3821), .B(N4001), .Y(N4049) );
  NOR2X1 gate1441 ( .A(N4005), .B(N4006), .Y(N4052) );
  NOR2X1 gate1442 ( .A(N4007), .B(N4008), .Y(N4055) );
  NOR2X1 gate1443 ( .A(N4009), .B(N4010), .Y(N4058) );
  NOR2X1 gate1444 ( .A(N4011), .B(N4012), .Y(N4061) );
  NOR2X1 gate1445 ( .A(N4013), .B(N4014), .Y(N4064) );
  NOR2X1 gate1446 ( .A(N4015), .B(N4016), .Y(N4067) );
  NOR2X1 gate1447 ( .A(N4017), .B(N4018), .Y(N4070) );
  NOR2X1 gate1448 ( .A(N4019), .B(N906), .Y(N4073) );
  NOR2X1 gate1449 ( .A(N3977), .B(N4022), .Y(N4077) );
  NOR2X1 gate1450 ( .A(N4022), .B(N954), .Y(N4078) );
  NOR2X1 gate1451 ( .A(N3868), .B(N4022), .Y(N4079) );
  NOR2X1 gate1452 ( .A(N4026), .B(N4027), .Y(N4082) );
  NOR2X1 gate1453 ( .A(N4031), .B(N4028), .Y(N4085) );
  NOR2X1 gate1454 ( .A(N3989), .B(N4034), .Y(N4089) );
  NOR2X1 gate1455 ( .A(N4034), .B(N3986), .Y(N4090) );
  NOR2X1 gate1456 ( .A(N4038), .B(N4039), .Y(N4091) );
  NOR2X1 gate1457 ( .A(N4040), .B(N1149), .Y(N4094) );
  NOR2X1 gate1458 ( .A(N3998), .B(N4043), .Y(N4098) );
  NOR2X1 gate1459 ( .A(N4043), .B(N1197), .Y(N4099) );
  NOR2X1 gate1460 ( .A(N3889), .B(N4043), .Y(N4100) );
  NOR2X1 gate1461 ( .A(N4047), .B(N4048), .Y(N4103) );
  NOR2X1 gate1462 ( .A(N1293), .B(N4049), .Y(N4106) );
  NOR2X1 gate1463 ( .A(N4052), .B(N570), .Y(N4110) );
  NOR2X1 gate1464 ( .A(N4055), .B(N618), .Y(N4114) );
  NOR2X1 gate1465 ( .A(N4058), .B(N666), .Y(N4118) );
  NOR2X1 gate1466 ( .A(N4061), .B(N714), .Y(N4122) );
  NOR2X1 gate1467 ( .A(N4064), .B(N762), .Y(N4126) );
  NOR2X1 gate1468 ( .A(N4067), .B(N810), .Y(N4130) );
  NOR2X1 gate1469 ( .A(N4070), .B(N858), .Y(N4134) );
  NOR2X1 gate1470 ( .A(N4019), .B(N4073), .Y(N4138) );
  NOR2X1 gate1471 ( .A(N4073), .B(N906), .Y(N4139) );
  NOR2X1 gate1472 ( .A(N3917), .B(N4073), .Y(N4140) );
  NOR2X1 gate1473 ( .A(N4077), .B(N4078), .Y(N4143) );
  NOR2X1 gate1474 ( .A(N4082), .B(N4079), .Y(N4146) );
  NOR2X1 gate1475 ( .A(N4031), .B(N4085), .Y(N4150) );
  NOR2X1 gate1476 ( .A(N4085), .B(N4028), .Y(N4151) );
  NOR2X1 gate1477 ( .A(N4089), .B(N4090), .Y(N4152) );
  NOR2X1 gate1478 ( .A(N4091), .B(N1101), .Y(N4155) );
  NOR2X1 gate1479 ( .A(N4040), .B(N4094), .Y(N4159) );
  NOR2X1 gate1480 ( .A(N4094), .B(N1149), .Y(N4160) );
  NOR2X1 gate1481 ( .A(N3938), .B(N4094), .Y(N4161) );
  NOR2X1 gate1482 ( .A(N4098), .B(N4099), .Y(N4164) );
  NOR2X1 gate1483 ( .A(N4103), .B(N4100), .Y(N4167) );
  NOR2X1 gate1484 ( .A(N1293), .B(N4106), .Y(N4171) );
  NOR2X1 gate1485 ( .A(N4106), .B(N4049), .Y(N4172) );
  NOR2X1 gate1486 ( .A(N4052), .B(N4110), .Y(N4173) );
  NOR2X1 gate1487 ( .A(N4110), .B(N570), .Y(N4174) );
  NOR2X1 gate1488 ( .A(N3947), .B(N4110), .Y(N4175) );
  NOR2X1 gate1489 ( .A(N4055), .B(N4114), .Y(N4178) );
  NOR2X1 gate1490 ( .A(N4114), .B(N618), .Y(N4179) );
  NOR2X1 gate1491 ( .A(N3951), .B(N4114), .Y(N4180) );
  NOR2X1 gate1492 ( .A(N4058), .B(N4118), .Y(N4183) );
  NOR2X1 gate1493 ( .A(N4118), .B(N666), .Y(N4184) );
  NOR2X1 gate1494 ( .A(N3955), .B(N4118), .Y(N4185) );
  NOR2X1 gate1495 ( .A(N4061), .B(N4122), .Y(N4188) );
  NOR2X1 gate1496 ( .A(N4122), .B(N714), .Y(N4189) );
  NOR2X1 gate1497 ( .A(N3959), .B(N4122), .Y(N4190) );
  NOR2X1 gate1498 ( .A(N4064), .B(N4126), .Y(N4193) );
  NOR2X1 gate1499 ( .A(N4126), .B(N762), .Y(N4194) );
  NOR2X1 gate1500 ( .A(N3963), .B(N4126), .Y(N4195) );
  NOR2X1 gate1501 ( .A(N4067), .B(N4130), .Y(N4198) );
  NOR2X1 gate1502 ( .A(N4130), .B(N810), .Y(N4199) );
  NOR2X1 gate1503 ( .A(N3967), .B(N4130), .Y(N4200) );
  NOR2X1 gate1504 ( .A(N4070), .B(N4134), .Y(N4203) );
  NOR2X1 gate1505 ( .A(N4134), .B(N858), .Y(N4204) );
  NOR2X1 gate1506 ( .A(N3971), .B(N4134), .Y(N4205) );
  NOR2X1 gate1507 ( .A(N4138), .B(N4139), .Y(N4208) );
  NOR2X1 gate1508 ( .A(N4143), .B(N4140), .Y(N4211) );
  NOR2X1 gate1509 ( .A(N4082), .B(N4146), .Y(N4215) );
  NOR2X1 gate1510 ( .A(N4146), .B(N4079), .Y(N4216) );
  NOR2X1 gate1511 ( .A(N4150), .B(N4151), .Y(N4217) );
  NOR2X1 gate1512 ( .A(N4152), .B(N1053), .Y(N4220) );
  NOR2X1 gate1513 ( .A(N4091), .B(N4155), .Y(N4224) );
  NOR2X1 gate1514 ( .A(N4155), .B(N1101), .Y(N4225) );
  NOR2X1 gate1515 ( .A(N3992), .B(N4155), .Y(N4226) );
  NOR2X1 gate1516 ( .A(N4159), .B(N4160), .Y(N4229) );
  NOR2X1 gate1517 ( .A(N4164), .B(N4161), .Y(N4232) );
  NOR2X1 gate1518 ( .A(N4103), .B(N4167), .Y(N4236) );
  NOR2X1 gate1519 ( .A(N4167), .B(N4100), .Y(N4237) );
  NOR2X1 gate1520 ( .A(N4171), .B(N4172), .Y(N4238) );
  NOR2X1 gate1521 ( .A(N4173), .B(N4174), .Y(N4241) );
  NOR2X1 gate1522 ( .A(N4178), .B(N4179), .Y(N4242) );
  NOR2X1 gate1523 ( .A(N4183), .B(N4184), .Y(N4245) );
  NOR2X1 gate1524 ( .A(N4188), .B(N4189), .Y(N4248) );
  NOR2X1 gate1525 ( .A(N4193), .B(N4194), .Y(N4251) );
  NOR2X1 gate1526 ( .A(N4198), .B(N4199), .Y(N4254) );
  NOR2X1 gate1527 ( .A(N4203), .B(N4204), .Y(N4257) );
  NOR2X1 gate1528 ( .A(N4208), .B(N4205), .Y(N4260) );
  NOR2X1 gate1529 ( .A(N4143), .B(N4211), .Y(N4264) );
  NOR2X1 gate1530 ( .A(N4211), .B(N4140), .Y(N4265) );
  NOR2X1 gate1531 ( .A(N4215), .B(N4216), .Y(N4266) );
  NOR2X1 gate1532 ( .A(N4217), .B(N1005), .Y(N4269) );
  NOR2X1 gate1533 ( .A(N4152), .B(N4220), .Y(N4273) );
  NOR2X1 gate1534 ( .A(N4220), .B(N1053), .Y(N4274) );
  NOR2X1 gate1535 ( .A(N4034), .B(N4220), .Y(N4275) );
  NOR2X1 gate1536 ( .A(N4224), .B(N4225), .Y(N4278) );
  NOR2X1 gate1537 ( .A(N4229), .B(N4226), .Y(N4281) );
  NOR2X1 gate1538 ( .A(N4164), .B(N4232), .Y(N4285) );
  NOR2X1 gate1539 ( .A(N4232), .B(N4161), .Y(N4286) );
  NOR2X1 gate1540 ( .A(N4236), .B(N4237), .Y(N4287) );
  NOR2X1 gate1541 ( .A(N4238), .B(N1248), .Y(N4290) );
  NOR2X1 gate1542 ( .A(N4242), .B(N4175), .Y(N4294) );
  NOR2X1 gate1543 ( .A(N4245), .B(N4180), .Y(N4298) );
  NOR2X1 gate1544 ( .A(N4248), .B(N4185), .Y(N4302) );
  NOR2X1 gate1545 ( .A(N4251), .B(N4190), .Y(N4306) );
  NOR2X1 gate1546 ( .A(N4254), .B(N4195), .Y(N4310) );
  NOR2X1 gate1547 ( .A(N4257), .B(N4200), .Y(N4314) );
  NOR2X1 gate1548 ( .A(N4208), .B(N4260), .Y(N4318) );
  NOR2X1 gate1549 ( .A(N4260), .B(N4205), .Y(N4319) );
  NOR2X1 gate1550 ( .A(N4264), .B(N4265), .Y(N4320) );
  NOR2X1 gate1551 ( .A(N4266), .B(N957), .Y(N4323) );
  NOR2X1 gate1552 ( .A(N4217), .B(N4269), .Y(N4327) );
  NOR2X1 gate1553 ( .A(N4269), .B(N1005), .Y(N4328) );
  NOR2X1 gate1554 ( .A(N4085), .B(N4269), .Y(N4329) );
  NOR2X1 gate1555 ( .A(N4273), .B(N4274), .Y(N4332) );
  NOR2X1 gate1556 ( .A(N4278), .B(N4275), .Y(N4335) );
  NOR2X1 gate1557 ( .A(N4229), .B(N4281), .Y(N4339) );
  NOR2X1 gate1558 ( .A(N4281), .B(N4226), .Y(N4340) );
  NOR2X1 gate1559 ( .A(N4285), .B(N4286), .Y(N4341) );
  NOR2X1 gate1560 ( .A(N4287), .B(N1200), .Y(N4344) );
  NOR2X1 gate1561 ( .A(N4238), .B(N4290), .Y(N4348) );
  NOR2X1 gate1562 ( .A(N4290), .B(N1248), .Y(N4349) );
  NOR2X1 gate1563 ( .A(N4106), .B(N4290), .Y(N4350) );
  NOR2X1 gate1564 ( .A(N4242), .B(N4294), .Y(N4353) );
  NOR2X1 gate1565 ( .A(N4294), .B(N4175), .Y(N4354) );
  NOR2X1 gate1566 ( .A(N4245), .B(N4298), .Y(N4355) );
  NOR2X1 gate1567 ( .A(N4298), .B(N4180), .Y(N4356) );
  NOR2X1 gate1568 ( .A(N4248), .B(N4302), .Y(N4357) );
  NOR2X1 gate1569 ( .A(N4302), .B(N4185), .Y(N4358) );
  NOR2X1 gate1570 ( .A(N4251), .B(N4306), .Y(N4359) );
  NOR2X1 gate1571 ( .A(N4306), .B(N4190), .Y(N4360) );
  NOR2X1 gate1572 ( .A(N4254), .B(N4310), .Y(N4361) );
  NOR2X1 gate1573 ( .A(N4310), .B(N4195), .Y(N4362) );
  NOR2X1 gate1574 ( .A(N4257), .B(N4314), .Y(N4363) );
  NOR2X1 gate1575 ( .A(N4314), .B(N4200), .Y(N4364) );
  NOR2X1 gate1576 ( .A(N4318), .B(N4319), .Y(N4365) );
  NOR2X1 gate1577 ( .A(N4320), .B(N909), .Y(N4368) );
  NOR2X1 gate1578 ( .A(N4266), .B(N4323), .Y(N4372) );
  NOR2X1 gate1579 ( .A(N4323), .B(N957), .Y(N4373) );
  NOR2X1 gate1580 ( .A(N4146), .B(N4323), .Y(N4374) );
  NOR2X1 gate1581 ( .A(N4327), .B(N4328), .Y(N4377) );
  NOR2X1 gate1582 ( .A(N4332), .B(N4329), .Y(N4380) );
  NOR2X1 gate1583 ( .A(N4278), .B(N4335), .Y(N4384) );
  NOR2X1 gate1584 ( .A(N4335), .B(N4275), .Y(N4385) );
  NOR2X1 gate1585 ( .A(N4339), .B(N4340), .Y(N4386) );
  NOR2X1 gate1586 ( .A(N4341), .B(N1152), .Y(N4389) );
  NOR2X1 gate1587 ( .A(N4287), .B(N4344), .Y(N4393) );
  NOR2X1 gate1588 ( .A(N4344), .B(N1200), .Y(N4394) );
  NOR2X1 gate1589 ( .A(N4167), .B(N4344), .Y(N4395) );
  NOR2X1 gate1590 ( .A(N4348), .B(N4349), .Y(N4398) );
  NOR2X1 gate1591 ( .A(N1296), .B(N4350), .Y(N4401) );
  NOR2X1 gate1592 ( .A(N4353), .B(N4354), .Y(N4405) );
  NOR2X1 gate1593 ( .A(N4355), .B(N4356), .Y(N4408) );
  NOR2X1 gate1594 ( .A(N4357), .B(N4358), .Y(N4411) );
  NOR2X1 gate1595 ( .A(N4359), .B(N4360), .Y(N4414) );
  NOR2X1 gate1596 ( .A(N4361), .B(N4362), .Y(N4417) );
  NOR2X1 gate1597 ( .A(N4363), .B(N4364), .Y(N4420) );
  NOR2X1 gate1598 ( .A(N4365), .B(N861), .Y(N4423) );
  NOR2X1 gate1599 ( .A(N4320), .B(N4368), .Y(N4427) );
  NOR2X1 gate1600 ( .A(N4368), .B(N909), .Y(N4428) );
  NOR2X1 gate1601 ( .A(N4211), .B(N4368), .Y(N4429) );
  NOR2X1 gate1602 ( .A(N4372), .B(N4373), .Y(N4432) );
  NOR2X1 gate1603 ( .A(N4377), .B(N4374), .Y(N4435) );
  NOR2X1 gate1604 ( .A(N4332), .B(N4380), .Y(N4439) );
  NOR2X1 gate1605 ( .A(N4380), .B(N4329), .Y(N4440) );
  NOR2X1 gate1606 ( .A(N4384), .B(N4385), .Y(N4441) );
  NOR2X1 gate1607 ( .A(N4386), .B(N1104), .Y(N4444) );
  NOR2X1 gate1608 ( .A(N4341), .B(N4389), .Y(N4448) );
  NOR2X1 gate1609 ( .A(N4389), .B(N1152), .Y(N4449) );
  NOR2X1 gate1610 ( .A(N4232), .B(N4389), .Y(N4450) );
  NOR2X1 gate1611 ( .A(N4393), .B(N4394), .Y(N4453) );
  NOR2X1 gate1612 ( .A(N4398), .B(N4395), .Y(N4456) );
  NOR2X1 gate1613 ( .A(N1296), .B(N4401), .Y(N4460) );
  NOR2X1 gate1614 ( .A(N4401), .B(N4350), .Y(N4461) );
  NOR2X1 gate1615 ( .A(N4405), .B(N573), .Y(N4462) );
  NOR2X1 gate1616 ( .A(N4408), .B(N621), .Y(N4466) );
  NOR2X1 gate1617 ( .A(N4411), .B(N669), .Y(N4470) );
  NOR2X1 gate1618 ( .A(N4414), .B(N717), .Y(N4474) );
  NOR2X1 gate1619 ( .A(N4417), .B(N765), .Y(N4478) );
  NOR2X1 gate1620 ( .A(N4420), .B(N813), .Y(N4482) );
  NOR2X1 gate1621 ( .A(N4365), .B(N4423), .Y(N4486) );
  NOR2X1 gate1622 ( .A(N4423), .B(N861), .Y(N4487) );
  NOR2X1 gate1623 ( .A(N4260), .B(N4423), .Y(N4488) );
  NOR2X1 gate1624 ( .A(N4427), .B(N4428), .Y(N4491) );
  NOR2X1 gate1625 ( .A(N4432), .B(N4429), .Y(N4494) );
  NOR2X1 gate1626 ( .A(N4377), .B(N4435), .Y(N4498) );
  NOR2X1 gate1627 ( .A(N4435), .B(N4374), .Y(N4499) );
  NOR2X1 gate1628 ( .A(N4439), .B(N4440), .Y(N4500) );
  NOR2X1 gate1629 ( .A(N4441), .B(N1056), .Y(N4503) );
  NOR2X1 gate1630 ( .A(N4386), .B(N4444), .Y(N4507) );
  NOR2X1 gate1631 ( .A(N4444), .B(N1104), .Y(N4508) );
  NOR2X1 gate1632 ( .A(N4281), .B(N4444), .Y(N4509) );
  NOR2X1 gate1633 ( .A(N4448), .B(N4449), .Y(N4512) );
  NOR2X1 gate1634 ( .A(N4453), .B(N4450), .Y(N4515) );
  NOR2X1 gate1635 ( .A(N4398), .B(N4456), .Y(N4519) );
  NOR2X1 gate1636 ( .A(N4456), .B(N4395), .Y(N4520) );
  NOR2X1 gate1637 ( .A(N4460), .B(N4461), .Y(N4521) );
  NOR2X1 gate1638 ( .A(N4405), .B(N4462), .Y(N4524) );
  NOR2X1 gate1639 ( .A(N4462), .B(N573), .Y(N4525) );
  NOR2X1 gate1640 ( .A(N4294), .B(N4462), .Y(N4526) );
  NOR2X1 gate1641 ( .A(N4408), .B(N4466), .Y(N4529) );
  NOR2X1 gate1642 ( .A(N4466), .B(N621), .Y(N4530) );
  NOR2X1 gate1643 ( .A(N4298), .B(N4466), .Y(N4531) );
  NOR2X1 gate1644 ( .A(N4411), .B(N4470), .Y(N4534) );
  NOR2X1 gate1645 ( .A(N4470), .B(N669), .Y(N4535) );
  NOR2X1 gate1646 ( .A(N4302), .B(N4470), .Y(N4536) );
  NOR2X1 gate1647 ( .A(N4414), .B(N4474), .Y(N4539) );
  NOR2X1 gate1648 ( .A(N4474), .B(N717), .Y(N4540) );
  NOR2X1 gate1649 ( .A(N4306), .B(N4474), .Y(N4541) );
  NOR2X1 gate1650 ( .A(N4417), .B(N4478), .Y(N4544) );
  NOR2X1 gate1651 ( .A(N4478), .B(N765), .Y(N4545) );
  NOR2X1 gate1652 ( .A(N4310), .B(N4478), .Y(N4546) );
  NOR2X1 gate1653 ( .A(N4420), .B(N4482), .Y(N4549) );
  NOR2X1 gate1654 ( .A(N4482), .B(N813), .Y(N4550) );
  NOR2X1 gate1655 ( .A(N4314), .B(N4482), .Y(N4551) );
  NOR2X1 gate1656 ( .A(N4486), .B(N4487), .Y(N4554) );
  NOR2X1 gate1657 ( .A(N4491), .B(N4488), .Y(N4557) );
  NOR2X1 gate1658 ( .A(N4432), .B(N4494), .Y(N4561) );
  NOR2X1 gate1659 ( .A(N4494), .B(N4429), .Y(N4562) );
  NOR2X1 gate1660 ( .A(N4498), .B(N4499), .Y(N4563) );
  NOR2X1 gate1661 ( .A(N4500), .B(N1008), .Y(N4566) );
  NOR2X1 gate1662 ( .A(N4441), .B(N4503), .Y(N4570) );
  NOR2X1 gate1663 ( .A(N4503), .B(N1056), .Y(N4571) );
  NOR2X1 gate1664 ( .A(N4335), .B(N4503), .Y(N4572) );
  NOR2X1 gate1665 ( .A(N4507), .B(N4508), .Y(N4575) );
  NOR2X1 gate1666 ( .A(N4512), .B(N4509), .Y(N4578) );
  NOR2X1 gate1667 ( .A(N4453), .B(N4515), .Y(N4582) );
  NOR2X1 gate1668 ( .A(N4515), .B(N4450), .Y(N4583) );
  NOR2X1 gate1669 ( .A(N4519), .B(N4520), .Y(N4584) );
  NOR2X1 gate1670 ( .A(N4521), .B(N1251), .Y(N4587) );
  NOR2X1 gate1671 ( .A(N4524), .B(N4525), .Y(N4591) );
  NOR2X1 gate1672 ( .A(N4529), .B(N4530), .Y(N4592) );
  NOR2X1 gate1673 ( .A(N4534), .B(N4535), .Y(N4595) );
  NOR2X1 gate1674 ( .A(N4539), .B(N4540), .Y(N4598) );
  NOR2X1 gate1675 ( .A(N4544), .B(N4545), .Y(N4601) );
  NOR2X1 gate1676 ( .A(N4549), .B(N4550), .Y(N4604) );
  NOR2X1 gate1677 ( .A(N4554), .B(N4551), .Y(N4607) );
  NOR2X1 gate1678 ( .A(N4491), .B(N4557), .Y(N4611) );
  NOR2X1 gate1679 ( .A(N4557), .B(N4488), .Y(N4612) );
  NOR2X1 gate1680 ( .A(N4561), .B(N4562), .Y(N4613) );
  NOR2X1 gate1681 ( .A(N4563), .B(N960), .Y(N4616) );
  NOR2X1 gate1682 ( .A(N4500), .B(N4566), .Y(N4620) );
  NOR2X1 gate1683 ( .A(N4566), .B(N1008), .Y(N4621) );
  NOR2X1 gate1684 ( .A(N4380), .B(N4566), .Y(N4622) );
  NOR2X1 gate1685 ( .A(N4570), .B(N4571), .Y(N4625) );
  NOR2X1 gate1686 ( .A(N4575), .B(N4572), .Y(N4628) );
  NOR2X1 gate1687 ( .A(N4512), .B(N4578), .Y(N4632) );
  NOR2X1 gate1688 ( .A(N4578), .B(N4509), .Y(N4633) );
  NOR2X1 gate1689 ( .A(N4582), .B(N4583), .Y(N4634) );
  NOR2X1 gate1690 ( .A(N4584), .B(N1203), .Y(N4637) );
  NOR2X1 gate1691 ( .A(N4521), .B(N4587), .Y(N4641) );
  NOR2X1 gate1692 ( .A(N4587), .B(N1251), .Y(N4642) );
  NOR2X1 gate1693 ( .A(N4401), .B(N4587), .Y(N4643) );
  NOR2X1 gate1694 ( .A(N4592), .B(N4526), .Y(N4646) );
  NOR2X1 gate1695 ( .A(N4595), .B(N4531), .Y(N4650) );
  NOR2X1 gate1696 ( .A(N4598), .B(N4536), .Y(N4654) );
  NOR2X1 gate1697 ( .A(N4601), .B(N4541), .Y(N4658) );
  NOR2X1 gate1698 ( .A(N4604), .B(N4546), .Y(N4662) );
  NOR2X1 gate1699 ( .A(N4554), .B(N4607), .Y(N4666) );
  NOR2X1 gate1700 ( .A(N4607), .B(N4551), .Y(N4667) );
  NOR2X1 gate1701 ( .A(N4611), .B(N4612), .Y(N4668) );
  NOR2X1 gate1702 ( .A(N4613), .B(N912), .Y(N4671) );
  NOR2X1 gate1703 ( .A(N4563), .B(N4616), .Y(N4675) );
  NOR2X1 gate1704 ( .A(N4616), .B(N960), .Y(N4676) );
  NOR2X1 gate1705 ( .A(N4435), .B(N4616), .Y(N4677) );
  NOR2X1 gate1706 ( .A(N4620), .B(N4621), .Y(N4680) );
  NOR2X1 gate1707 ( .A(N4625), .B(N4622), .Y(N4683) );
  NOR2X1 gate1708 ( .A(N4575), .B(N4628), .Y(N4687) );
  NOR2X1 gate1709 ( .A(N4628), .B(N4572), .Y(N4688) );
  NOR2X1 gate1710 ( .A(N4632), .B(N4633), .Y(N4689) );
  NOR2X1 gate1711 ( .A(N4634), .B(N1155), .Y(N4692) );
  NOR2X1 gate1712 ( .A(N4584), .B(N4637), .Y(N4696) );
  NOR2X1 gate1713 ( .A(N4637), .B(N1203), .Y(N4697) );
  NOR2X1 gate1714 ( .A(N4456), .B(N4637), .Y(N4698) );
  NOR2X1 gate1715 ( .A(N4641), .B(N4642), .Y(N4701) );
  NOR2X1 gate1716 ( .A(N1299), .B(N4643), .Y(N4704) );
  NOR2X1 gate1717 ( .A(N4592), .B(N4646), .Y(N4708) );
  NOR2X1 gate1718 ( .A(N4646), .B(N4526), .Y(N4709) );
  NOR2X1 gate1719 ( .A(N4595), .B(N4650), .Y(N4710) );
  NOR2X1 gate1720 ( .A(N4650), .B(N4531), .Y(N4711) );
  NOR2X1 gate1721 ( .A(N4598), .B(N4654), .Y(N4712) );
  NOR2X1 gate1722 ( .A(N4654), .B(N4536), .Y(N4713) );
  NOR2X1 gate1723 ( .A(N4601), .B(N4658), .Y(N4714) );
  NOR2X1 gate1724 ( .A(N4658), .B(N4541), .Y(N4715) );
  NOR2X1 gate1725 ( .A(N4604), .B(N4662), .Y(N4716) );
  NOR2X1 gate1726 ( .A(N4662), .B(N4546), .Y(N4717) );
  NOR2X1 gate1727 ( .A(N4666), .B(N4667), .Y(N4718) );
  NOR2X1 gate1728 ( .A(N4668), .B(N864), .Y(N4721) );
  NOR2X1 gate1729 ( .A(N4613), .B(N4671), .Y(N4725) );
  NOR2X1 gate1730 ( .A(N4671), .B(N912), .Y(N4726) );
  NOR2X1 gate1731 ( .A(N4494), .B(N4671), .Y(N4727) );
  NOR2X1 gate1732 ( .A(N4675), .B(N4676), .Y(N4730) );
  NOR2X1 gate1733 ( .A(N4680), .B(N4677), .Y(N4733) );
  NOR2X1 gate1734 ( .A(N4625), .B(N4683), .Y(N4737) );
  NOR2X1 gate1735 ( .A(N4683), .B(N4622), .Y(N4738) );
  NOR2X1 gate1736 ( .A(N4687), .B(N4688), .Y(N4739) );
  NOR2X1 gate1737 ( .A(N4689), .B(N1107), .Y(N4742) );
  NOR2X1 gate1738 ( .A(N4634), .B(N4692), .Y(N4746) );
  NOR2X1 gate1739 ( .A(N4692), .B(N1155), .Y(N4747) );
  NOR2X1 gate1740 ( .A(N4515), .B(N4692), .Y(N4748) );
  NOR2X1 gate1741 ( .A(N4696), .B(N4697), .Y(N4751) );
  NOR2X1 gate1742 ( .A(N4701), .B(N4698), .Y(N4754) );
  NOR2X1 gate1743 ( .A(N1299), .B(N4704), .Y(N4758) );
  NOR2X1 gate1744 ( .A(N4704), .B(N4643), .Y(N4759) );
  NOR2X1 gate1745 ( .A(N4708), .B(N4709), .Y(N4760) );
  NOR2X1 gate1746 ( .A(N4710), .B(N4711), .Y(N4763) );
  NOR2X1 gate1747 ( .A(N4712), .B(N4713), .Y(N4766) );
  NOR2X1 gate1748 ( .A(N4714), .B(N4715), .Y(N4769) );
  NOR2X1 gate1749 ( .A(N4716), .B(N4717), .Y(N4772) );
  NOR2X1 gate1750 ( .A(N4718), .B(N816), .Y(N4775) );
  NOR2X1 gate1751 ( .A(N4668), .B(N4721), .Y(N4779) );
  NOR2X1 gate1752 ( .A(N4721), .B(N864), .Y(N4780) );
  NOR2X1 gate1753 ( .A(N4557), .B(N4721), .Y(N4781) );
  NOR2X1 gate1754 ( .A(N4725), .B(N4726), .Y(N4784) );
  NOR2X1 gate1755 ( .A(N4730), .B(N4727), .Y(N4787) );
  NOR2X1 gate1756 ( .A(N4680), .B(N4733), .Y(N4791) );
  NOR2X1 gate1757 ( .A(N4733), .B(N4677), .Y(N4792) );
  NOR2X1 gate1758 ( .A(N4737), .B(N4738), .Y(N4793) );
  NOR2X1 gate1759 ( .A(N4739), .B(N1059), .Y(N4796) );
  NOR2X1 gate1760 ( .A(N4689), .B(N4742), .Y(N4800) );
  NOR2X1 gate1761 ( .A(N4742), .B(N1107), .Y(N4801) );
  NOR2X1 gate1762 ( .A(N4578), .B(N4742), .Y(N4802) );
  NOR2X1 gate1763 ( .A(N4746), .B(N4747), .Y(N4805) );
  NOR2X1 gate1764 ( .A(N4751), .B(N4748), .Y(N4808) );
  NOR2X1 gate1765 ( .A(N4701), .B(N4754), .Y(N4812) );
  NOR2X1 gate1766 ( .A(N4754), .B(N4698), .Y(N4813) );
  NOR2X1 gate1767 ( .A(N4758), .B(N4759), .Y(N4814) );
  NOR2X1 gate1768 ( .A(N4760), .B(N576), .Y(N4817) );
  NOR2X1 gate1769 ( .A(N4763), .B(N624), .Y(N4821) );
  NOR2X1 gate1770 ( .A(N4766), .B(N672), .Y(N4825) );
  NOR2X1 gate1771 ( .A(N4769), .B(N720), .Y(N4829) );
  NOR2X1 gate1772 ( .A(N4772), .B(N768), .Y(N4833) );
  NOR2X1 gate1773 ( .A(N4718), .B(N4775), .Y(N4837) );
  NOR2X1 gate1774 ( .A(N4775), .B(N816), .Y(N4838) );
  NOR2X1 gate1775 ( .A(N4607), .B(N4775), .Y(N4839) );
  NOR2X1 gate1776 ( .A(N4779), .B(N4780), .Y(N4842) );
  NOR2X1 gate1777 ( .A(N4784), .B(N4781), .Y(N4845) );
  NOR2X1 gate1778 ( .A(N4730), .B(N4787), .Y(N4849) );
  NOR2X1 gate1779 ( .A(N4787), .B(N4727), .Y(N4850) );
  NOR2X1 gate1780 ( .A(N4791), .B(N4792), .Y(N4851) );
  NOR2X1 gate1781 ( .A(N4793), .B(N1011), .Y(N4854) );
  NOR2X1 gate1782 ( .A(N4739), .B(N4796), .Y(N4858) );
  NOR2X1 gate1783 ( .A(N4796), .B(N1059), .Y(N4859) );
  NOR2X1 gate1784 ( .A(N4628), .B(N4796), .Y(N4860) );
  NOR2X1 gate1785 ( .A(N4800), .B(N4801), .Y(N4863) );
  NOR2X1 gate1786 ( .A(N4805), .B(N4802), .Y(N4866) );
  NOR2X1 gate1787 ( .A(N4751), .B(N4808), .Y(N4870) );
  NOR2X1 gate1788 ( .A(N4808), .B(N4748), .Y(N4871) );
  NOR2X1 gate1789 ( .A(N4812), .B(N4813), .Y(N4872) );
  NOR2X1 gate1790 ( .A(N4814), .B(N1254), .Y(N4875) );
  NOR2X1 gate1791 ( .A(N4760), .B(N4817), .Y(N4879) );
  NOR2X1 gate1792 ( .A(N4817), .B(N576), .Y(N4880) );
  NOR2X1 gate1793 ( .A(N4646), .B(N4817), .Y(N4881) );
  NOR2X1 gate1794 ( .A(N4763), .B(N4821), .Y(N4884) );
  NOR2X1 gate1795 ( .A(N4821), .B(N624), .Y(N4885) );
  NOR2X1 gate1796 ( .A(N4650), .B(N4821), .Y(N4886) );
  NOR2X1 gate1797 ( .A(N4766), .B(N4825), .Y(N4889) );
  NOR2X1 gate1798 ( .A(N4825), .B(N672), .Y(N4890) );
  NOR2X1 gate1799 ( .A(N4654), .B(N4825), .Y(N4891) );
  NOR2X1 gate1800 ( .A(N4769), .B(N4829), .Y(N4894) );
  NOR2X1 gate1801 ( .A(N4829), .B(N720), .Y(N4895) );
  NOR2X1 gate1802 ( .A(N4658), .B(N4829), .Y(N4896) );
  NOR2X1 gate1803 ( .A(N4772), .B(N4833), .Y(N4899) );
  NOR2X1 gate1804 ( .A(N4833), .B(N768), .Y(N4900) );
  NOR2X1 gate1805 ( .A(N4662), .B(N4833), .Y(N4901) );
  NOR2X1 gate1806 ( .A(N4837), .B(N4838), .Y(N4904) );
  NOR2X1 gate1807 ( .A(N4842), .B(N4839), .Y(N4907) );
  NOR2X1 gate1808 ( .A(N4784), .B(N4845), .Y(N4911) );
  NOR2X1 gate1809 ( .A(N4845), .B(N4781), .Y(N4912) );
  NOR2X1 gate1810 ( .A(N4849), .B(N4850), .Y(N4913) );
  NOR2X1 gate1811 ( .A(N4851), .B(N963), .Y(N4916) );
  NOR2X1 gate1812 ( .A(N4793), .B(N4854), .Y(N4920) );
  NOR2X1 gate1813 ( .A(N4854), .B(N1011), .Y(N4921) );
  NOR2X1 gate1814 ( .A(N4683), .B(N4854), .Y(N4922) );
  NOR2X1 gate1815 ( .A(N4858), .B(N4859), .Y(N4925) );
  NOR2X1 gate1816 ( .A(N4863), .B(N4860), .Y(N4928) );
  NOR2X1 gate1817 ( .A(N4805), .B(N4866), .Y(N4932) );
  NOR2X1 gate1818 ( .A(N4866), .B(N4802), .Y(N4933) );
  NOR2X1 gate1819 ( .A(N4870), .B(N4871), .Y(N4934) );
  NOR2X1 gate1820 ( .A(N4872), .B(N1206), .Y(N4937) );
  NOR2X1 gate1821 ( .A(N4814), .B(N4875), .Y(N4941) );
  NOR2X1 gate1822 ( .A(N4875), .B(N1254), .Y(N4942) );
  NOR2X1 gate1823 ( .A(N4704), .B(N4875), .Y(N4943) );
  NOR2X1 gate1824 ( .A(N4879), .B(N4880), .Y(N4946) );
  NOR2X1 gate1825 ( .A(N4884), .B(N4885), .Y(N4947) );
  NOR2X1 gate1826 ( .A(N4889), .B(N4890), .Y(N4950) );
  NOR2X1 gate1827 ( .A(N4894), .B(N4895), .Y(N4953) );
  NOR2X1 gate1828 ( .A(N4899), .B(N4900), .Y(N4956) );
  NOR2X1 gate1829 ( .A(N4904), .B(N4901), .Y(N4959) );
  NOR2X1 gate1830 ( .A(N4842), .B(N4907), .Y(N4963) );
  NOR2X1 gate1831 ( .A(N4907), .B(N4839), .Y(N4964) );
  NOR2X1 gate1832 ( .A(N4911), .B(N4912), .Y(N4965) );
  NOR2X1 gate1833 ( .A(N4913), .B(N915), .Y(N4968) );
  NOR2X1 gate1834 ( .A(N4851), .B(N4916), .Y(N4972) );
  NOR2X1 gate1835 ( .A(N4916), .B(N963), .Y(N4973) );
  NOR2X1 gate1836 ( .A(N4733), .B(N4916), .Y(N4974) );
  NOR2X1 gate1837 ( .A(N4920), .B(N4921), .Y(N4977) );
  NOR2X1 gate1838 ( .A(N4925), .B(N4922), .Y(N4980) );
  NOR2X1 gate1839 ( .A(N4863), .B(N4928), .Y(N4984) );
  NOR2X1 gate1840 ( .A(N4928), .B(N4860), .Y(N4985) );
  NOR2X1 gate1841 ( .A(N4932), .B(N4933), .Y(N4986) );
  NOR2X1 gate1842 ( .A(N4934), .B(N1158), .Y(N4989) );
  NOR2X1 gate1843 ( .A(N4872), .B(N4937), .Y(N4993) );
  NOR2X1 gate1844 ( .A(N4937), .B(N1206), .Y(N4994) );
  NOR2X1 gate1845 ( .A(N4754), .B(N4937), .Y(N4995) );
  NOR2X1 gate1846 ( .A(N4941), .B(N4942), .Y(N4998) );
  NOR2X1 gate1847 ( .A(N1302), .B(N4943), .Y(N5001) );
  NOR2X1 gate1848 ( .A(N4947), .B(N4881), .Y(N5005) );
  NOR2X1 gate1849 ( .A(N4950), .B(N4886), .Y(N5009) );
  NOR2X1 gate1850 ( .A(N4953), .B(N4891), .Y(N5013) );
  NOR2X1 gate1851 ( .A(N4956), .B(N4896), .Y(N5017) );
  NOR2X1 gate1852 ( .A(N4904), .B(N4959), .Y(N5021) );
  NOR2X1 gate1853 ( .A(N4959), .B(N4901), .Y(N5022) );
  NOR2X1 gate1854 ( .A(N4963), .B(N4964), .Y(N5023) );
  NOR2X1 gate1855 ( .A(N4965), .B(N867), .Y(N5026) );
  NOR2X1 gate1856 ( .A(N4913), .B(N4968), .Y(N5030) );
  NOR2X1 gate1857 ( .A(N4968), .B(N915), .Y(N5031) );
  NOR2X1 gate1858 ( .A(N4787), .B(N4968), .Y(N5032) );
  NOR2X1 gate1859 ( .A(N4972), .B(N4973), .Y(N5035) );
  NOR2X1 gate1860 ( .A(N4977), .B(N4974), .Y(N5038) );
  NOR2X1 gate1861 ( .A(N4925), .B(N4980), .Y(N5042) );
  NOR2X1 gate1862 ( .A(N4980), .B(N4922), .Y(N5043) );
  NOR2X1 gate1863 ( .A(N4984), .B(N4985), .Y(N5044) );
  NOR2X1 gate1864 ( .A(N4986), .B(N1110), .Y(N5047) );
  NOR2X1 gate1865 ( .A(N4934), .B(N4989), .Y(N5051) );
  NOR2X1 gate1866 ( .A(N4989), .B(N1158), .Y(N5052) );
  NOR2X1 gate1867 ( .A(N4808), .B(N4989), .Y(N5053) );
  NOR2X1 gate1868 ( .A(N4993), .B(N4994), .Y(N5056) );
  NOR2X1 gate1869 ( .A(N4998), .B(N4995), .Y(N5059) );
  NOR2X1 gate1870 ( .A(N1302), .B(N5001), .Y(N5063) );
  NOR2X1 gate1871 ( .A(N5001), .B(N4943), .Y(N5064) );
  NOR2X1 gate1872 ( .A(N4947), .B(N5005), .Y(N5065) );
  NOR2X1 gate1873 ( .A(N5005), .B(N4881), .Y(N5066) );
  NOR2X1 gate1874 ( .A(N4950), .B(N5009), .Y(N5067) );
  NOR2X1 gate1875 ( .A(N5009), .B(N4886), .Y(N5068) );
  NOR2X1 gate1876 ( .A(N4953), .B(N5013), .Y(N5069) );
  NOR2X1 gate1877 ( .A(N5013), .B(N4891), .Y(N5070) );
  NOR2X1 gate1878 ( .A(N4956), .B(N5017), .Y(N5071) );
  NOR2X1 gate1879 ( .A(N5017), .B(N4896), .Y(N5072) );
  NOR2X1 gate1880 ( .A(N5021), .B(N5022), .Y(N5073) );
  NOR2X1 gate1881 ( .A(N5023), .B(N819), .Y(N5076) );
  NOR2X1 gate1882 ( .A(N4965), .B(N5026), .Y(N5080) );
  NOR2X1 gate1883 ( .A(N5026), .B(N867), .Y(N5081) );
  NOR2X1 gate1884 ( .A(N4845), .B(N5026), .Y(N5082) );
  NOR2X1 gate1885 ( .A(N5030), .B(N5031), .Y(N5085) );
  NOR2X1 gate1886 ( .A(N5035), .B(N5032), .Y(N5088) );
  NOR2X1 gate1887 ( .A(N4977), .B(N5038), .Y(N5092) );
  NOR2X1 gate1888 ( .A(N5038), .B(N4974), .Y(N5093) );
  NOR2X1 gate1889 ( .A(N5042), .B(N5043), .Y(N5094) );
  NOR2X1 gate1890 ( .A(N5044), .B(N1062), .Y(N5097) );
  NOR2X1 gate1891 ( .A(N4986), .B(N5047), .Y(N5101) );
  NOR2X1 gate1892 ( .A(N5047), .B(N1110), .Y(N5102) );
  NOR2X1 gate1893 ( .A(N4866), .B(N5047), .Y(N5103) );
  NOR2X1 gate1894 ( .A(N5051), .B(N5052), .Y(N5106) );
  NOR2X1 gate1895 ( .A(N5056), .B(N5053), .Y(N5109) );
  NOR2X1 gate1896 ( .A(N4998), .B(N5059), .Y(N5113) );
  NOR2X1 gate1897 ( .A(N5059), .B(N4995), .Y(N5114) );
  NOR2X1 gate1898 ( .A(N5063), .B(N5064), .Y(N5115) );
  NOR2X1 gate1899 ( .A(N5065), .B(N5066), .Y(N5118) );
  NOR2X1 gate1900 ( .A(N5067), .B(N5068), .Y(N5121) );
  NOR2X1 gate1901 ( .A(N5069), .B(N5070), .Y(N5124) );
  NOR2X1 gate1902 ( .A(N5071), .B(N5072), .Y(N5127) );
  NOR2X1 gate1903 ( .A(N5073), .B(N771), .Y(N5130) );
  NOR2X1 gate1904 ( .A(N5023), .B(N5076), .Y(N5134) );
  NOR2X1 gate1905 ( .A(N5076), .B(N819), .Y(N5135) );
  NOR2X1 gate1906 ( .A(N4907), .B(N5076), .Y(N5136) );
  NOR2X1 gate1907 ( .A(N5080), .B(N5081), .Y(N5139) );
  NOR2X1 gate1908 ( .A(N5085), .B(N5082), .Y(N5142) );
  NOR2X1 gate1909 ( .A(N5035), .B(N5088), .Y(N5146) );
  NOR2X1 gate1910 ( .A(N5088), .B(N5032), .Y(N5147) );
  NOR2X1 gate1911 ( .A(N5092), .B(N5093), .Y(N5148) );
  NOR2X1 gate1912 ( .A(N5094), .B(N1014), .Y(N5151) );
  NOR2X1 gate1913 ( .A(N5044), .B(N5097), .Y(N5155) );
  NOR2X1 gate1914 ( .A(N5097), .B(N1062), .Y(N5156) );
  NOR2X1 gate1915 ( .A(N4928), .B(N5097), .Y(N5157) );
  NOR2X1 gate1916 ( .A(N5101), .B(N5102), .Y(N5160) );
  NOR2X1 gate1917 ( .A(N5106), .B(N5103), .Y(N5163) );
  NOR2X1 gate1918 ( .A(N5056), .B(N5109), .Y(N5167) );
  NOR2X1 gate1919 ( .A(N5109), .B(N5053), .Y(N5168) );
  NOR2X1 gate1920 ( .A(N5113), .B(N5114), .Y(N5169) );
  NOR2X1 gate1921 ( .A(N5115), .B(N1257), .Y(N5172) );
  NOR2X1 gate1922 ( .A(N5118), .B(N579), .Y(N5176) );
  NOR2X1 gate1923 ( .A(N5121), .B(N627), .Y(N5180) );
  NOR2X1 gate1924 ( .A(N5124), .B(N675), .Y(N5184) );
  NOR2X1 gate1925 ( .A(N5127), .B(N723), .Y(N5188) );
  NOR2X1 gate1926 ( .A(N5073), .B(N5130), .Y(N5192) );
  NOR2X1 gate1927 ( .A(N5130), .B(N771), .Y(N5193) );
  NOR2X1 gate1928 ( .A(N4959), .B(N5130), .Y(N5194) );
  NOR2X1 gate1929 ( .A(N5134), .B(N5135), .Y(N5197) );
  NOR2X1 gate1930 ( .A(N5139), .B(N5136), .Y(N5200) );
  NOR2X1 gate1931 ( .A(N5085), .B(N5142), .Y(N5204) );
  NOR2X1 gate1932 ( .A(N5142), .B(N5082), .Y(N5205) );
  NOR2X1 gate1933 ( .A(N5146), .B(N5147), .Y(N5206) );
  NOR2X1 gate1934 ( .A(N5148), .B(N966), .Y(N5209) );
  NOR2X1 gate1935 ( .A(N5094), .B(N5151), .Y(N5213) );
  NOR2X1 gate1936 ( .A(N5151), .B(N1014), .Y(N5214) );
  NOR2X1 gate1937 ( .A(N4980), .B(N5151), .Y(N5215) );
  NOR2X1 gate1938 ( .A(N5155), .B(N5156), .Y(N5218) );
  NOR2X1 gate1939 ( .A(N5160), .B(N5157), .Y(N5221) );
  NOR2X1 gate1940 ( .A(N5106), .B(N5163), .Y(N5225) );
  NOR2X1 gate1941 ( .A(N5163), .B(N5103), .Y(N5226) );
  NOR2X1 gate1942 ( .A(N5167), .B(N5168), .Y(N5227) );
  NOR2X1 gate1943 ( .A(N5169), .B(N1209), .Y(N5230) );
  NOR2X1 gate1944 ( .A(N5115), .B(N5172), .Y(N5234) );
  NOR2X1 gate1945 ( .A(N5172), .B(N1257), .Y(N5235) );
  NOR2X1 gate1946 ( .A(N5001), .B(N5172), .Y(N5236) );
  NOR2X1 gate1947 ( .A(N5118), .B(N5176), .Y(N5239) );
  NOR2X1 gate1948 ( .A(N5176), .B(N579), .Y(N5240) );
  NOR2X1 gate1949 ( .A(N5005), .B(N5176), .Y(N5241) );
  NOR2X1 gate1950 ( .A(N5121), .B(N5180), .Y(N5244) );
  NOR2X1 gate1951 ( .A(N5180), .B(N627), .Y(N5245) );
  NOR2X1 gate1952 ( .A(N5009), .B(N5180), .Y(N5246) );
  NOR2X1 gate1953 ( .A(N5124), .B(N5184), .Y(N5249) );
  NOR2X1 gate1954 ( .A(N5184), .B(N675), .Y(N5250) );
  NOR2X1 gate1955 ( .A(N5013), .B(N5184), .Y(N5251) );
  NOR2X1 gate1956 ( .A(N5127), .B(N5188), .Y(N5254) );
  NOR2X1 gate1957 ( .A(N5188), .B(N723), .Y(N5255) );
  NOR2X1 gate1958 ( .A(N5017), .B(N5188), .Y(N5256) );
  NOR2X1 gate1959 ( .A(N5192), .B(N5193), .Y(N5259) );
  NOR2X1 gate1960 ( .A(N5197), .B(N5194), .Y(N5262) );
  NOR2X1 gate1961 ( .A(N5139), .B(N5200), .Y(N5266) );
  NOR2X1 gate1962 ( .A(N5200), .B(N5136), .Y(N5267) );
  NOR2X1 gate1963 ( .A(N5204), .B(N5205), .Y(N5268) );
  NOR2X1 gate1964 ( .A(N5206), .B(N918), .Y(N5271) );
  NOR2X1 gate1965 ( .A(N5148), .B(N5209), .Y(N5275) );
  NOR2X1 gate1966 ( .A(N5209), .B(N966), .Y(N5276) );
  NOR2X1 gate1967 ( .A(N5038), .B(N5209), .Y(N5277) );
  NOR2X1 gate1968 ( .A(N5213), .B(N5214), .Y(N5280) );
  NOR2X1 gate1969 ( .A(N5218), .B(N5215), .Y(N5283) );
  NOR2X1 gate1970 ( .A(N5160), .B(N5221), .Y(N5287) );
  NOR2X1 gate1971 ( .A(N5221), .B(N5157), .Y(N5288) );
  NOR2X1 gate1972 ( .A(N5225), .B(N5226), .Y(N5289) );
  NOR2X1 gate1973 ( .A(N5227), .B(N1161), .Y(N5292) );
  NOR2X1 gate1974 ( .A(N5169), .B(N5230), .Y(N5296) );
  NOR2X1 gate1975 ( .A(N5230), .B(N1209), .Y(N5297) );
  NOR2X1 gate1976 ( .A(N5059), .B(N5230), .Y(N5298) );
  NOR2X1 gate1977 ( .A(N5234), .B(N5235), .Y(N5301) );
  NOR2X1 gate1978 ( .A(N1305), .B(N5236), .Y(N5304) );
  NOR2X1 gate1979 ( .A(N5239), .B(N5240), .Y(N5308) );
  NOR2X1 gate1980 ( .A(N5244), .B(N5245), .Y(N5309) );
  NOR2X1 gate1981 ( .A(N5249), .B(N5250), .Y(N5312) );
  NOR2X1 gate1982 ( .A(N5254), .B(N5255), .Y(N5315) );
  NOR2X1 gate1983 ( .A(N5259), .B(N5256), .Y(N5318) );
  NOR2X1 gate1984 ( .A(N5197), .B(N5262), .Y(N5322) );
  NOR2X1 gate1985 ( .A(N5262), .B(N5194), .Y(N5323) );
  NOR2X1 gate1986 ( .A(N5266), .B(N5267), .Y(N5324) );
  NOR2X1 gate1987 ( .A(N5268), .B(N870), .Y(N5327) );
  NOR2X1 gate1988 ( .A(N5206), .B(N5271), .Y(N5331) );
  NOR2X1 gate1989 ( .A(N5271), .B(N918), .Y(N5332) );
  NOR2X1 gate1990 ( .A(N5088), .B(N5271), .Y(N5333) );
  NOR2X1 gate1991 ( .A(N5275), .B(N5276), .Y(N5336) );
  NOR2X1 gate1992 ( .A(N5280), .B(N5277), .Y(N5339) );
  NOR2X1 gate1993 ( .A(N5218), .B(N5283), .Y(N5343) );
  NOR2X1 gate1994 ( .A(N5283), .B(N5215), .Y(N5344) );
  NOR2X1 gate1995 ( .A(N5287), .B(N5288), .Y(N5345) );
  NOR2X1 gate1996 ( .A(N5289), .B(N1113), .Y(N5348) );
  NOR2X1 gate1997 ( .A(N5227), .B(N5292), .Y(N5352) );
  NOR2X1 gate1998 ( .A(N5292), .B(N1161), .Y(N5353) );
  NOR2X1 gate1999 ( .A(N5109), .B(N5292), .Y(N5354) );
  NOR2X1 gate2000 ( .A(N5296), .B(N5297), .Y(N5357) );
  NOR2X1 gate2001 ( .A(N5301), .B(N5298), .Y(N5360) );
  NOR2X1 gate2002 ( .A(N1305), .B(N5304), .Y(N5364) );
  NOR2X1 gate2003 ( .A(N5304), .B(N5236), .Y(N5365) );
  NOR2X1 gate2004 ( .A(N5309), .B(N5241), .Y(N5366) );
  NOR2X1 gate2005 ( .A(N5312), .B(N5246), .Y(N5370) );
  NOR2X1 gate2006 ( .A(N5315), .B(N5251), .Y(N5374) );
  NOR2X1 gate2007 ( .A(N5259), .B(N5318), .Y(N5378) );
  NOR2X1 gate2008 ( .A(N5318), .B(N5256), .Y(N5379) );
  NOR2X1 gate2009 ( .A(N5322), .B(N5323), .Y(N5380) );
  NOR2X1 gate2010 ( .A(N5324), .B(N822), .Y(N5383) );
  NOR2X1 gate2011 ( .A(N5268), .B(N5327), .Y(N5387) );
  NOR2X1 gate2012 ( .A(N5327), .B(N870), .Y(N5388) );
  NOR2X1 gate2013 ( .A(N5142), .B(N5327), .Y(N5389) );
  NOR2X1 gate2014 ( .A(N5331), .B(N5332), .Y(N5392) );
  NOR2X1 gate2015 ( .A(N5336), .B(N5333), .Y(N5395) );
  NOR2X1 gate2016 ( .A(N5280), .B(N5339), .Y(N5399) );
  NOR2X1 gate2017 ( .A(N5339), .B(N5277), .Y(N5400) );
  NOR2X1 gate2018 ( .A(N5343), .B(N5344), .Y(N5401) );
  NOR2X1 gate2019 ( .A(N5345), .B(N1065), .Y(N5404) );
  NOR2X1 gate2020 ( .A(N5289), .B(N5348), .Y(N5408) );
  NOR2X1 gate2021 ( .A(N5348), .B(N1113), .Y(N5409) );
  NOR2X1 gate2022 ( .A(N5163), .B(N5348), .Y(N5410) );
  NOR2X1 gate2023 ( .A(N5352), .B(N5353), .Y(N5413) );
  NOR2X1 gate2024 ( .A(N5357), .B(N5354), .Y(N5416) );
  NOR2X1 gate2025 ( .A(N5301), .B(N5360), .Y(N5420) );
  NOR2X1 gate2026 ( .A(N5360), .B(N5298), .Y(N5421) );
  NOR2X1 gate2027 ( .A(N5364), .B(N5365), .Y(N5422) );
  NOR2X1 gate2028 ( .A(N5309), .B(N5366), .Y(N5425) );
  NOR2X1 gate2029 ( .A(N5366), .B(N5241), .Y(N5426) );
  NOR2X1 gate2030 ( .A(N5312), .B(N5370), .Y(N5427) );
  NOR2X1 gate2031 ( .A(N5370), .B(N5246), .Y(N5428) );
  NOR2X1 gate2032 ( .A(N5315), .B(N5374), .Y(N5429) );
  NOR2X1 gate2033 ( .A(N5374), .B(N5251), .Y(N5430) );
  NOR2X1 gate2034 ( .A(N5378), .B(N5379), .Y(N5431) );
  NOR2X1 gate2035 ( .A(N5380), .B(N774), .Y(N5434) );
  NOR2X1 gate2036 ( .A(N5324), .B(N5383), .Y(N5438) );
  NOR2X1 gate2037 ( .A(N5383), .B(N822), .Y(N5439) );
  NOR2X1 gate2038 ( .A(N5200), .B(N5383), .Y(N5440) );
  NOR2X1 gate2039 ( .A(N5387), .B(N5388), .Y(N5443) );
  NOR2X1 gate2040 ( .A(N5392), .B(N5389), .Y(N5446) );
  NOR2X1 gate2041 ( .A(N5336), .B(N5395), .Y(N5450) );
  NOR2X1 gate2042 ( .A(N5395), .B(N5333), .Y(N5451) );
  NOR2X1 gate2043 ( .A(N5399), .B(N5400), .Y(N5452) );
  NOR2X1 gate2044 ( .A(N5401), .B(N1017), .Y(N5455) );
  NOR2X1 gate2045 ( .A(N5345), .B(N5404), .Y(N5459) );
  NOR2X1 gate2046 ( .A(N5404), .B(N1065), .Y(N5460) );
  NOR2X1 gate2047 ( .A(N5221), .B(N5404), .Y(N5461) );
  NOR2X1 gate2048 ( .A(N5408), .B(N5409), .Y(N5464) );
  NOR2X1 gate2049 ( .A(N5413), .B(N5410), .Y(N5467) );
  NOR2X1 gate2050 ( .A(N5357), .B(N5416), .Y(N5471) );
  NOR2X1 gate2051 ( .A(N5416), .B(N5354), .Y(N5472) );
  NOR2X1 gate2052 ( .A(N5420), .B(N5421), .Y(N5473) );
  NOR2X1 gate2053 ( .A(N5422), .B(N1260), .Y(N5476) );
  NOR2X1 gate2054 ( .A(N5425), .B(N5426), .Y(N5480) );
  NOR2X1 gate2055 ( .A(N5427), .B(N5428), .Y(N5483) );
  NOR2X1 gate2056 ( .A(N5429), .B(N5430), .Y(N5486) );
  NOR2X1 gate2057 ( .A(N5431), .B(N726), .Y(N5489) );
  NOR2X1 gate2058 ( .A(N5380), .B(N5434), .Y(N5493) );
  NOR2X1 gate2059 ( .A(N5434), .B(N774), .Y(N5494) );
  NOR2X1 gate2060 ( .A(N5262), .B(N5434), .Y(N5495) );
  NOR2X1 gate2061 ( .A(N5438), .B(N5439), .Y(N5498) );
  NOR2X1 gate2062 ( .A(N5443), .B(N5440), .Y(N5501) );
  NOR2X1 gate2063 ( .A(N5392), .B(N5446), .Y(N5505) );
  NOR2X1 gate2064 ( .A(N5446), .B(N5389), .Y(N5506) );
  NOR2X1 gate2065 ( .A(N5450), .B(N5451), .Y(N5507) );
  NOR2X1 gate2066 ( .A(N5452), .B(N969), .Y(N5510) );
  NOR2X1 gate2067 ( .A(N5401), .B(N5455), .Y(N5514) );
  NOR2X1 gate2068 ( .A(N5455), .B(N1017), .Y(N5515) );
  NOR2X1 gate2069 ( .A(N5283), .B(N5455), .Y(N5516) );
  NOR2X1 gate2070 ( .A(N5459), .B(N5460), .Y(N5519) );
  NOR2X1 gate2071 ( .A(N5464), .B(N5461), .Y(N5522) );
  NOR2X1 gate2072 ( .A(N5413), .B(N5467), .Y(N5526) );
  NOR2X1 gate2073 ( .A(N5467), .B(N5410), .Y(N5527) );
  NOR2X1 gate2074 ( .A(N5471), .B(N5472), .Y(N5528) );
  NOR2X1 gate2075 ( .A(N5473), .B(N1212), .Y(N5531) );
  NOR2X1 gate2076 ( .A(N5422), .B(N5476), .Y(N5535) );
  NOR2X1 gate2077 ( .A(N5476), .B(N1260), .Y(N5536) );
  NOR2X1 gate2078 ( .A(N5304), .B(N5476), .Y(N5537) );
  NOR2X1 gate2079 ( .A(N5480), .B(N582), .Y(N5540) );
  NOR2X1 gate2080 ( .A(N5483), .B(N630), .Y(N5544) );
  NOR2X1 gate2081 ( .A(N5486), .B(N678), .Y(N5548) );
  NOR2X1 gate2082 ( .A(N5431), .B(N5489), .Y(N5552) );
  NOR2X1 gate2083 ( .A(N5489), .B(N726), .Y(N5553) );
  NOR2X1 gate2084 ( .A(N5318), .B(N5489), .Y(N5554) );
  NOR2X1 gate2085 ( .A(N5493), .B(N5494), .Y(N5557) );
  NOR2X1 gate2086 ( .A(N5498), .B(N5495), .Y(N5560) );
  NOR2X1 gate2087 ( .A(N5443), .B(N5501), .Y(N5564) );
  NOR2X1 gate2088 ( .A(N5501), .B(N5440), .Y(N5565) );
  NOR2X1 gate2089 ( .A(N5505), .B(N5506), .Y(N5566) );
  NOR2X1 gate2090 ( .A(N5507), .B(N921), .Y(N5569) );
  NOR2X1 gate2091 ( .A(N5452), .B(N5510), .Y(N5573) );
  NOR2X1 gate2092 ( .A(N5510), .B(N969), .Y(N5574) );
  NOR2X1 gate2093 ( .A(N5339), .B(N5510), .Y(N5575) );
  NOR2X1 gate2094 ( .A(N5514), .B(N5515), .Y(N5578) );
  NOR2X1 gate2095 ( .A(N5519), .B(N5516), .Y(N5581) );
  NOR2X1 gate2096 ( .A(N5464), .B(N5522), .Y(N5585) );
  NOR2X1 gate2097 ( .A(N5522), .B(N5461), .Y(N5586) );
  NOR2X1 gate2098 ( .A(N5526), .B(N5527), .Y(N5587) );
  NOR2X1 gate2099 ( .A(N5528), .B(N1164), .Y(N5590) );
  NOR2X1 gate2100 ( .A(N5473), .B(N5531), .Y(N5594) );
  NOR2X1 gate2101 ( .A(N5531), .B(N1212), .Y(N5595) );
  NOR2X1 gate2102 ( .A(N5360), .B(N5531), .Y(N5596) );
  NOR2X1 gate2103 ( .A(N5535), .B(N5536), .Y(N5599) );
  NOR2X1 gate2104 ( .A(N1308), .B(N5537), .Y(N5602) );
  NOR2X1 gate2105 ( .A(N5480), .B(N5540), .Y(N5606) );
  NOR2X1 gate2106 ( .A(N5540), .B(N582), .Y(N5607) );
  NOR2X1 gate2107 ( .A(N5366), .B(N5540), .Y(N5608) );
  NOR2X1 gate2108 ( .A(N5483), .B(N5544), .Y(N5611) );
  NOR2X1 gate2109 ( .A(N5544), .B(N630), .Y(N5612) );
  NOR2X1 gate2110 ( .A(N5370), .B(N5544), .Y(N5613) );
  NOR2X1 gate2111 ( .A(N5486), .B(N5548), .Y(N5616) );
  NOR2X1 gate2112 ( .A(N5548), .B(N678), .Y(N5617) );
  NOR2X1 gate2113 ( .A(N5374), .B(N5548), .Y(N5618) );
  NOR2X1 gate2114 ( .A(N5552), .B(N5553), .Y(N5621) );
  NOR2X1 gate2115 ( .A(N5557), .B(N5554), .Y(N5624) );
  NOR2X1 gate2116 ( .A(N5498), .B(N5560), .Y(N5628) );
  NOR2X1 gate2117 ( .A(N5560), .B(N5495), .Y(N5629) );
  NOR2X1 gate2118 ( .A(N5564), .B(N5565), .Y(N5630) );
  NOR2X1 gate2119 ( .A(N5566), .B(N873), .Y(N5633) );
  NOR2X1 gate2120 ( .A(N5507), .B(N5569), .Y(N5637) );
  NOR2X1 gate2121 ( .A(N5569), .B(N921), .Y(N5638) );
  NOR2X1 gate2122 ( .A(N5395), .B(N5569), .Y(N5639) );
  NOR2X1 gate2123 ( .A(N5573), .B(N5574), .Y(N5642) );
  NOR2X1 gate2124 ( .A(N5578), .B(N5575), .Y(N5645) );
  NOR2X1 gate2125 ( .A(N5519), .B(N5581), .Y(N5649) );
  NOR2X1 gate2126 ( .A(N5581), .B(N5516), .Y(N5650) );
  NOR2X1 gate2127 ( .A(N5585), .B(N5586), .Y(N5651) );
  NOR2X1 gate2128 ( .A(N5587), .B(N1116), .Y(N5654) );
  NOR2X1 gate2129 ( .A(N5528), .B(N5590), .Y(N5658) );
  NOR2X1 gate2130 ( .A(N5590), .B(N1164), .Y(N5659) );
  NOR2X1 gate2131 ( .A(N5416), .B(N5590), .Y(N5660) );
  NOR2X1 gate2132 ( .A(N5594), .B(N5595), .Y(N5663) );
  NOR2X1 gate2133 ( .A(N5599), .B(N5596), .Y(N5666) );
  NOR2X1 gate2134 ( .A(N1308), .B(N5602), .Y(N5670) );
  NOR2X1 gate2135 ( .A(N5602), .B(N5537), .Y(N5671) );
  NOR2X1 gate2136 ( .A(N5606), .B(N5607), .Y(N5672) );
  NOR2X1 gate2137 ( .A(N5611), .B(N5612), .Y(N5673) );
  NOR2X1 gate2138 ( .A(N5616), .B(N5617), .Y(N5676) );
  NOR2X1 gate2139 ( .A(N5621), .B(N5618), .Y(N5679) );
  NOR2X1 gate2140 ( .A(N5557), .B(N5624), .Y(N5683) );
  NOR2X1 gate2141 ( .A(N5624), .B(N5554), .Y(N5684) );
  NOR2X1 gate2142 ( .A(N5628), .B(N5629), .Y(N5685) );
  NOR2X1 gate2143 ( .A(N5630), .B(N825), .Y(N5688) );
  NOR2X1 gate2144 ( .A(N5566), .B(N5633), .Y(N5692) );
  NOR2X1 gate2145 ( .A(N5633), .B(N873), .Y(N5693) );
  NOR2X1 gate2146 ( .A(N5446), .B(N5633), .Y(N5694) );
  NOR2X1 gate2147 ( .A(N5637), .B(N5638), .Y(N5697) );
  NOR2X1 gate2148 ( .A(N5642), .B(N5639), .Y(N5700) );
  NOR2X1 gate2149 ( .A(N5578), .B(N5645), .Y(N5704) );
  NOR2X1 gate2150 ( .A(N5645), .B(N5575), .Y(N5705) );
  NOR2X1 gate2151 ( .A(N5649), .B(N5650), .Y(N5706) );
  NOR2X1 gate2152 ( .A(N5651), .B(N1068), .Y(N5709) );
  NOR2X1 gate2153 ( .A(N5587), .B(N5654), .Y(N5713) );
  NOR2X1 gate2154 ( .A(N5654), .B(N1116), .Y(N5714) );
  NOR2X1 gate2155 ( .A(N5467), .B(N5654), .Y(N5715) );
  NOR2X1 gate2156 ( .A(N5658), .B(N5659), .Y(N5718) );
  NOR2X1 gate2157 ( .A(N5663), .B(N5660), .Y(N5721) );
  NOR2X1 gate2158 ( .A(N5599), .B(N5666), .Y(N5725) );
  NOR2X1 gate2159 ( .A(N5666), .B(N5596), .Y(N5726) );
  NOR2X1 gate2160 ( .A(N5670), .B(N5671), .Y(N5727) );
  NOR2X1 gate2161 ( .A(N5673), .B(N5608), .Y(N5730) );
  NOR2X1 gate2162 ( .A(N5676), .B(N5613), .Y(N5734) );
  NOR2X1 gate2163 ( .A(N5621), .B(N5679), .Y(N5738) );
  NOR2X1 gate2164 ( .A(N5679), .B(N5618), .Y(N5739) );
  NOR2X1 gate2165 ( .A(N5683), .B(N5684), .Y(N5740) );
  NOR2X1 gate2166 ( .A(N5685), .B(N777), .Y(N5743) );
  NOR2X1 gate2167 ( .A(N5630), .B(N5688), .Y(N5747) );
  NOR2X1 gate2168 ( .A(N5688), .B(N825), .Y(N5748) );
  NOR2X1 gate2169 ( .A(N5501), .B(N5688), .Y(N5749) );
  NOR2X1 gate2170 ( .A(N5692), .B(N5693), .Y(N5752) );
  NOR2X1 gate2171 ( .A(N5697), .B(N5694), .Y(N5755) );
  NOR2X1 gate2172 ( .A(N5642), .B(N5700), .Y(N5759) );
  NOR2X1 gate2173 ( .A(N5700), .B(N5639), .Y(N5760) );
  NOR2X1 gate2174 ( .A(N5704), .B(N5705), .Y(N5761) );
  NOR2X1 gate2175 ( .A(N5706), .B(N1020), .Y(N5764) );
  NOR2X1 gate2176 ( .A(N5651), .B(N5709), .Y(N5768) );
  NOR2X1 gate2177 ( .A(N5709), .B(N1068), .Y(N5769) );
  NOR2X1 gate2178 ( .A(N5522), .B(N5709), .Y(N5770) );
  NOR2X1 gate2179 ( .A(N5713), .B(N5714), .Y(N5773) );
  NOR2X1 gate2180 ( .A(N5718), .B(N5715), .Y(N5776) );
  NOR2X1 gate2181 ( .A(N5663), .B(N5721), .Y(N5780) );
  NOR2X1 gate2182 ( .A(N5721), .B(N5660), .Y(N5781) );
  NOR2X1 gate2183 ( .A(N5725), .B(N5726), .Y(N5782) );
  NOR2X1 gate2184 ( .A(N5673), .B(N5730), .Y(N5785) );
  NOR2X1 gate2185 ( .A(N5730), .B(N5608), .Y(N5786) );
  NOR2X1 gate2186 ( .A(N5676), .B(N5734), .Y(N5787) );
  NOR2X1 gate2187 ( .A(N5734), .B(N5613), .Y(N5788) );
  NOR2X1 gate2188 ( .A(N5738), .B(N5739), .Y(N5789) );
  NOR2X1 gate2189 ( .A(N5740), .B(N729), .Y(N5792) );
  NOR2X1 gate2190 ( .A(N5685), .B(N5743), .Y(N5796) );
  NOR2X1 gate2191 ( .A(N5743), .B(N777), .Y(N5797) );
  NOR2X1 gate2192 ( .A(N5560), .B(N5743), .Y(N5798) );
  NOR2X1 gate2193 ( .A(N5747), .B(N5748), .Y(N5801) );
  NOR2X1 gate2194 ( .A(N5752), .B(N5749), .Y(N5804) );
  NOR2X1 gate2195 ( .A(N5697), .B(N5755), .Y(N5808) );
  NOR2X1 gate2196 ( .A(N5755), .B(N5694), .Y(N5809) );
  NOR2X1 gate2197 ( .A(N5759), .B(N5760), .Y(N5810) );
  NOR2X1 gate2198 ( .A(N5761), .B(N972), .Y(N5813) );
  NOR2X1 gate2199 ( .A(N5706), .B(N5764), .Y(N5817) );
  NOR2X1 gate2200 ( .A(N5764), .B(N1020), .Y(N5818) );
  NOR2X1 gate2201 ( .A(N5581), .B(N5764), .Y(N5819) );
  NOR2X1 gate2202 ( .A(N5768), .B(N5769), .Y(N5822) );
  NOR2X1 gate2203 ( .A(N5773), .B(N5770), .Y(N5825) );
  NOR2X1 gate2204 ( .A(N5718), .B(N5776), .Y(N5829) );
  NOR2X1 gate2205 ( .A(N5776), .B(N5715), .Y(N5830) );
  NOR2X1 gate2206 ( .A(N5780), .B(N5781), .Y(N5831) );
  NOR2X1 gate2207 ( .A(N5785), .B(N5786), .Y(N5834) );
  NOR2X1 gate2208 ( .A(N5787), .B(N5788), .Y(N5837) );
  NOR2X1 gate2209 ( .A(N5789), .B(N681), .Y(N5840) );
  NOR2X1 gate2210 ( .A(N5740), .B(N5792), .Y(N5844) );
  NOR2X1 gate2211 ( .A(N5792), .B(N729), .Y(N5845) );
  NOR2X1 gate2212 ( .A(N5624), .B(N5792), .Y(N5846) );
  NOR2X1 gate2213 ( .A(N5796), .B(N5797), .Y(N5849) );
  NOR2X1 gate2214 ( .A(N5801), .B(N5798), .Y(N5852) );
  NOR2X1 gate2215 ( .A(N5752), .B(N5804), .Y(N5856) );
  NOR2X1 gate2216 ( .A(N5804), .B(N5749), .Y(N5857) );
  NOR2X1 gate2217 ( .A(N5808), .B(N5809), .Y(N5858) );
  NOR2X1 gate2218 ( .A(N5810), .B(N924), .Y(N5861) );
  NOR2X1 gate2219 ( .A(N5761), .B(N5813), .Y(N5865) );
  NOR2X1 gate2220 ( .A(N5813), .B(N972), .Y(N5866) );
  NOR2X1 gate2221 ( .A(N5645), .B(N5813), .Y(N5867) );
  NOR2X1 gate2222 ( .A(N5817), .B(N5818), .Y(N5870) );
  NOR2X1 gate2223 ( .A(N5822), .B(N5819), .Y(N5873) );
  NOR2X1 gate2224 ( .A(N5773), .B(N5825), .Y(N5877) );
  NOR2X1 gate2225 ( .A(N5825), .B(N5770), .Y(N5878) );
  NOR2X1 gate2226 ( .A(N5829), .B(N5830), .Y(N5879) );
  NOR2X1 gate2227 ( .A(N5834), .B(N585), .Y(N5882) );
  NOR2X1 gate2228 ( .A(N5837), .B(N633), .Y(N5886) );
  NOR2X1 gate2229 ( .A(N5789), .B(N5840), .Y(N5890) );
  NOR2X1 gate2230 ( .A(N5840), .B(N681), .Y(N5891) );
  NOR2X1 gate2231 ( .A(N5679), .B(N5840), .Y(N5892) );
  NOR2X1 gate2232 ( .A(N5844), .B(N5845), .Y(N5895) );
  NOR2X1 gate2233 ( .A(N5849), .B(N5846), .Y(N5898) );
  NOR2X1 gate2234 ( .A(N5801), .B(N5852), .Y(N5902) );
  NOR2X1 gate2235 ( .A(N5852), .B(N5798), .Y(N5903) );
  NOR2X1 gate2236 ( .A(N5856), .B(N5857), .Y(N5904) );
  NOR2X1 gate2237 ( .A(N5858), .B(N876), .Y(N5907) );
  NOR2X1 gate2238 ( .A(N5810), .B(N5861), .Y(N5911) );
  NOR2X1 gate2239 ( .A(N5861), .B(N924), .Y(N5912) );
  NOR2X1 gate2240 ( .A(N5700), .B(N5861), .Y(N5913) );
  NOR2X1 gate2241 ( .A(N5865), .B(N5866), .Y(N5916) );
  NOR2X1 gate2242 ( .A(N5870), .B(N5867), .Y(N5919) );
  NOR2X1 gate2243 ( .A(N5822), .B(N5873), .Y(N5923) );
  NOR2X1 gate2244 ( .A(N5873), .B(N5819), .Y(N5924) );
  NOR2X1 gate2245 ( .A(N5877), .B(N5878), .Y(N5925) );
  NOR2X1 gate2246 ( .A(N5834), .B(N5882), .Y(N5928) );
  NOR2X1 gate2247 ( .A(N5882), .B(N585), .Y(N5929) );
  NOR2X1 gate2248 ( .A(N5730), .B(N5882), .Y(N5930) );
  NOR2X1 gate2249 ( .A(N5837), .B(N5886), .Y(N5933) );
  NOR2X1 gate2250 ( .A(N5886), .B(N633), .Y(N5934) );
  NOR2X1 gate2251 ( .A(N5734), .B(N5886), .Y(N5935) );
  NOR2X1 gate2252 ( .A(N5890), .B(N5891), .Y(N5938) );
  NOR2X1 gate2253 ( .A(N5895), .B(N5892), .Y(N5941) );
  NOR2X1 gate2254 ( .A(N5849), .B(N5898), .Y(N5945) );
  NOR2X1 gate2255 ( .A(N5898), .B(N5846), .Y(N5946) );
  NOR2X1 gate2256 ( .A(N5902), .B(N5903), .Y(N5947) );
  NOR2X1 gate2257 ( .A(N5904), .B(N828), .Y(N5950) );
  NOR2X1 gate2258 ( .A(N5858), .B(N5907), .Y(N5954) );
  NOR2X1 gate2259 ( .A(N5907), .B(N876), .Y(N5955) );
  NOR2X1 gate2260 ( .A(N5755), .B(N5907), .Y(N5956) );
  NOR2X1 gate2261 ( .A(N5911), .B(N5912), .Y(N5959) );
  NOR2X1 gate2262 ( .A(N5916), .B(N5913), .Y(N5962) );
  NOR2X1 gate2263 ( .A(N5870), .B(N5919), .Y(N5966) );
  NOR2X1 gate2264 ( .A(N5919), .B(N5867), .Y(N5967) );
  NOR2X1 gate2265 ( .A(N5923), .B(N5924), .Y(N5968) );
  NOR2X1 gate2266 ( .A(N5928), .B(N5929), .Y(N5971) );
  NOR2X1 gate2267 ( .A(N5933), .B(N5934), .Y(N5972) );
  NOR2X1 gate2268 ( .A(N5938), .B(N5935), .Y(N5975) );
  NOR2X1 gate2269 ( .A(N5895), .B(N5941), .Y(N5979) );
  NOR2X1 gate2270 ( .A(N5941), .B(N5892), .Y(N5980) );
  NOR2X1 gate2271 ( .A(N5945), .B(N5946), .Y(N5981) );
  NOR2X1 gate2272 ( .A(N5947), .B(N780), .Y(N5984) );
  NOR2X1 gate2273 ( .A(N5904), .B(N5950), .Y(N5988) );
  NOR2X1 gate2274 ( .A(N5950), .B(N828), .Y(N5989) );
  NOR2X1 gate2275 ( .A(N5804), .B(N5950), .Y(N5990) );
  NOR2X1 gate2276 ( .A(N5954), .B(N5955), .Y(N5993) );
  NOR2X1 gate2277 ( .A(N5959), .B(N5956), .Y(N5996) );
  NOR2X1 gate2278 ( .A(N5916), .B(N5962), .Y(N6000) );
  NOR2X1 gate2279 ( .A(N5962), .B(N5913), .Y(N6001) );
  NOR2X1 gate2280 ( .A(N5966), .B(N5967), .Y(N6002) );
  NOR2X1 gate2281 ( .A(N5972), .B(N5930), .Y(N6005) );
  NOR2X1 gate2282 ( .A(N5938), .B(N5975), .Y(N6009) );
  NOR2X1 gate2283 ( .A(N5975), .B(N5935), .Y(N6010) );
  NOR2X1 gate2284 ( .A(N5979), .B(N5980), .Y(N6011) );
  NOR2X1 gate2285 ( .A(N5981), .B(N732), .Y(N6014) );
  NOR2X1 gate2286 ( .A(N5947), .B(N5984), .Y(N6018) );
  NOR2X1 gate2287 ( .A(N5984), .B(N780), .Y(N6019) );
  NOR2X1 gate2288 ( .A(N5852), .B(N5984), .Y(N6020) );
  NOR2X1 gate2289 ( .A(N5988), .B(N5989), .Y(N6023) );
  NOR2X1 gate2290 ( .A(N5993), .B(N5990), .Y(N6026) );
  NOR2X1 gate2291 ( .A(N5959), .B(N5996), .Y(N6030) );
  NOR2X1 gate2292 ( .A(N5996), .B(N5956), .Y(N6031) );
  NOR2X1 gate2293 ( .A(N6000), .B(N6001), .Y(N6032) );
  NOR2X1 gate2294 ( .A(N5972), .B(N6005), .Y(N6035) );
  NOR2X1 gate2295 ( .A(N6005), .B(N5930), .Y(N6036) );
  NOR2X1 gate2296 ( .A(N6009), .B(N6010), .Y(N6037) );
  NOR2X1 gate2297 ( .A(N6011), .B(N684), .Y(N6040) );
  NOR2X1 gate2298 ( .A(N5981), .B(N6014), .Y(N6044) );
  NOR2X1 gate2299 ( .A(N6014), .B(N732), .Y(N6045) );
  NOR2X1 gate2300 ( .A(N5898), .B(N6014), .Y(N6046) );
  NOR2X1 gate2301 ( .A(N6018), .B(N6019), .Y(N6049) );
  NOR2X1 gate2302 ( .A(N6023), .B(N6020), .Y(N6052) );
  NOR2X1 gate2303 ( .A(N5993), .B(N6026), .Y(N6056) );
  NOR2X1 gate2304 ( .A(N6026), .B(N5990), .Y(N6057) );
  NOR2X1 gate2305 ( .A(N6030), .B(N6031), .Y(N6058) );
  NOR2X1 gate2306 ( .A(N6035), .B(N6036), .Y(N6061) );
  NOR2X1 gate2307 ( .A(N6037), .B(N636), .Y(N6064) );
  NOR2X1 gate2308 ( .A(N6011), .B(N6040), .Y(N6068) );
  NOR2X1 gate2309 ( .A(N6040), .B(N684), .Y(N6069) );
  NOR2X1 gate2310 ( .A(N5941), .B(N6040), .Y(N6070) );
  NOR2X1 gate2311 ( .A(N6044), .B(N6045), .Y(N6073) );
  NOR2X1 gate2312 ( .A(N6049), .B(N6046), .Y(N6076) );
  NOR2X1 gate2313 ( .A(N6023), .B(N6052), .Y(N6080) );
  NOR2X1 gate2314 ( .A(N6052), .B(N6020), .Y(N6081) );
  NOR2X1 gate2315 ( .A(N6056), .B(N6057), .Y(N6082) );
  NOR2X1 gate2316 ( .A(N6061), .B(N588), .Y(N6085) );
  NOR2X1 gate2317 ( .A(N6037), .B(N6064), .Y(N6089) );
  NOR2X1 gate2318 ( .A(N6064), .B(N636), .Y(N6090) );
  NOR2X1 gate2319 ( .A(N5975), .B(N6064), .Y(N6091) );
  NOR2X1 gate2320 ( .A(N6068), .B(N6069), .Y(N6094) );
  NOR2X1 gate2321 ( .A(N6073), .B(N6070), .Y(N6097) );
  NOR2X1 gate2322 ( .A(N6049), .B(N6076), .Y(N6101) );
  NOR2X1 gate2323 ( .A(N6076), .B(N6046), .Y(N6102) );
  NOR2X1 gate2324 ( .A(N6080), .B(N6081), .Y(N6103) );
  NOR2X1 gate2325 ( .A(N6061), .B(N6085), .Y(N6106) );
  NOR2X1 gate2326 ( .A(N6085), .B(N588), .Y(N6107) );
  NOR2X1 gate2327 ( .A(N6005), .B(N6085), .Y(N6108) );
  NOR2X1 gate2328 ( .A(N6089), .B(N6090), .Y(N6111) );
  NOR2X1 gate2329 ( .A(N6094), .B(N6091), .Y(N6114) );
  NOR2X1 gate2330 ( .A(N6073), .B(N6097), .Y(N6118) );
  NOR2X1 gate2331 ( .A(N6097), .B(N6070), .Y(N6119) );
  NOR2X1 gate2332 ( .A(N6101), .B(N6102), .Y(N6120) );
  NOR2X1 gate2333 ( .A(N6106), .B(N6107), .Y(N6123) );
  NOR2X1 gate2334 ( .A(N6111), .B(N6108), .Y(N6124) );
  NOR2X1 gate2335 ( .A(N6094), .B(N6114), .Y(N6128) );
  NOR2X1 gate2336 ( .A(N6114), .B(N6091), .Y(N6129) );
  NOR2X1 gate2337 ( .A(N6118), .B(N6119), .Y(N6130) );
  NOR2X1 gate2338 ( .A(N6111), .B(N6124), .Y(N6133) );
  NOR2X1 gate2339 ( .A(N6124), .B(N6108), .Y(N6134) );
  NOR2X1 gate2340 ( .A(N6128), .B(N6129), .Y(N6135) );
  NOR2X1 gate2341 ( .A(N6133), .B(N6134), .Y(N6138) );
  INVX1 gate2342 ( .A(N6138), .Y(N6141) );
  NOR2X1 gate2343 ( .A(N6138), .B(N6141), .Y(N6145) );
  INVX1 gate2344 ( .A(N6141), .Y(N6146) );
  NOR2X1 gate2345 ( .A(N6124), .B(N6141), .Y(N6147) );
  NOR2X1 gate2346 ( .A(N6145), .B(N6146), .Y(N6150) );
  NOR2X1 gate2347 ( .A(N6135), .B(N6147), .Y(N6151) );
  NOR2X1 gate2348 ( .A(N6135), .B(N6151), .Y(N6155) );
  NOR2X1 gate2349 ( .A(N6151), .B(N6147), .Y(N6156) );
  NOR2X1 gate2350 ( .A(N6114), .B(N6151), .Y(N6157) );
  NOR2X1 gate2351 ( .A(N6155), .B(N6156), .Y(N6160) );
  NOR2X1 gate2352 ( .A(N6130), .B(N6157), .Y(N6161) );
  NOR2X1 gate2353 ( .A(N6130), .B(N6161), .Y(N6165) );
  NOR2X1 gate2354 ( .A(N6161), .B(N6157), .Y(N6166) );
  NOR2X1 gate2355 ( .A(N6097), .B(N6161), .Y(N6167) );
  NOR2X1 gate2356 ( .A(N6165), .B(N6166), .Y(N6170) );
  NOR2X1 gate2357 ( .A(N6120), .B(N6167), .Y(N6171) );
  NOR2X1 gate2358 ( .A(N6120), .B(N6171), .Y(N6175) );
  NOR2X1 gate2359 ( .A(N6171), .B(N6167), .Y(N6176) );
  NOR2X1 gate2360 ( .A(N6076), .B(N6171), .Y(N6177) );
  NOR2X1 gate2361 ( .A(N6175), .B(N6176), .Y(N6180) );
  NOR2X1 gate2362 ( .A(N6103), .B(N6177), .Y(N6181) );
  NOR2X1 gate2363 ( .A(N6103), .B(N6181), .Y(N6185) );
  NOR2X1 gate2364 ( .A(N6181), .B(N6177), .Y(N6186) );
  NOR2X1 gate2365 ( .A(N6052), .B(N6181), .Y(N6187) );
  NOR2X1 gate2366 ( .A(N6185), .B(N6186), .Y(N6190) );
  NOR2X1 gate2367 ( .A(N6082), .B(N6187), .Y(N6191) );
  NOR2X1 gate2368 ( .A(N6082), .B(N6191), .Y(N6195) );
  NOR2X1 gate2369 ( .A(N6191), .B(N6187), .Y(N6196) );
  NOR2X1 gate2370 ( .A(N6026), .B(N6191), .Y(N6197) );
  NOR2X1 gate2371 ( .A(N6195), .B(N6196), .Y(N6200) );
  NOR2X1 gate2372 ( .A(N6058), .B(N6197), .Y(N6201) );
  NOR2X1 gate2373 ( .A(N6058), .B(N6201), .Y(N6205) );
  NOR2X1 gate2374 ( .A(N6201), .B(N6197), .Y(N6206) );
  NOR2X1 gate2375 ( .A(N5996), .B(N6201), .Y(N6207) );
  NOR2X1 gate2376 ( .A(N6205), .B(N6206), .Y(N6210) );
  NOR2X1 gate2377 ( .A(N6032), .B(N6207), .Y(N6211) );
  NOR2X1 gate2378 ( .A(N6032), .B(N6211), .Y(N6215) );
  NOR2X1 gate2379 ( .A(N6211), .B(N6207), .Y(N6216) );
  NOR2X1 gate2380 ( .A(N5962), .B(N6211), .Y(N6217) );
  NOR2X1 gate2381 ( .A(N6215), .B(N6216), .Y(N6220) );
  NOR2X1 gate2382 ( .A(N6002), .B(N6217), .Y(N6221) );
  NOR2X1 gate2383 ( .A(N6002), .B(N6221), .Y(N6225) );
  NOR2X1 gate2384 ( .A(N6221), .B(N6217), .Y(N6226) );
  NOR2X1 gate2385 ( .A(N5919), .B(N6221), .Y(N6227) );
  NOR2X1 gate2386 ( .A(N6225), .B(N6226), .Y(N6230) );
  NOR2X1 gate2387 ( .A(N5968), .B(N6227), .Y(N6231) );
  NOR2X1 gate2388 ( .A(N5968), .B(N6231), .Y(N6235) );
  NOR2X1 gate2389 ( .A(N6231), .B(N6227), .Y(N6236) );
  NOR2X1 gate2390 ( .A(N5873), .B(N6231), .Y(N6237) );
  NOR2X1 gate2391 ( .A(N6235), .B(N6236), .Y(N6240) );
  NOR2X1 gate2392 ( .A(N5925), .B(N6237), .Y(N6241) );
  NOR2X1 gate2393 ( .A(N5925), .B(N6241), .Y(N6245) );
  NOR2X1 gate2394 ( .A(N6241), .B(N6237), .Y(N6246) );
  NOR2X1 gate2395 ( .A(N5825), .B(N6241), .Y(N6247) );
  NOR2X1 gate2396 ( .A(N6245), .B(N6246), .Y(N6250) );
  NOR2X1 gate2397 ( .A(N5879), .B(N6247), .Y(N6251) );
  NOR2X1 gate2398 ( .A(N5879), .B(N6251), .Y(N6255) );
  NOR2X1 gate2399 ( .A(N6251), .B(N6247), .Y(N6256) );
  NOR2X1 gate2400 ( .A(N5776), .B(N6251), .Y(N6257) );
  NOR2X1 gate2401 ( .A(N6255), .B(N6256), .Y(N6260) );
  NOR2X1 gate2402 ( .A(N5831), .B(N6257), .Y(N6261) );
  NOR2X1 gate2403 ( .A(N5831), .B(N6261), .Y(N6265) );
  NOR2X1 gate2404 ( .A(N6261), .B(N6257), .Y(N6266) );
  NOR2X1 gate2405 ( .A(N5721), .B(N6261), .Y(N6267) );
  NOR2X1 gate2406 ( .A(N6265), .B(N6266), .Y(N6270) );
  NOR2X1 gate2407 ( .A(N5782), .B(N6267), .Y(N6271) );
  NOR2X1 gate2408 ( .A(N5782), .B(N6271), .Y(N6275) );
  NOR2X1 gate2409 ( .A(N6271), .B(N6267), .Y(N6276) );
  NOR2X1 gate2410 ( .A(N5666), .B(N6271), .Y(N6277) );
  NOR2X1 gate2411 ( .A(N6275), .B(N6276), .Y(N6280) );
  NOR2X1 gate2412 ( .A(N5727), .B(N6277), .Y(N6281) );
  NOR2X1 gate2413 ( .A(N5727), .B(N6281), .Y(N6285) );
  NOR2X1 gate2414 ( .A(N6281), .B(N6277), .Y(N6286) );
  NOR2X1 gate2415 ( .A(N5602), .B(N6281), .Y(N6287) );
  NOR2X1 gate2416 ( .A(N6285), .B(N6286), .Y(N6288) );
endmodule



module c2670_synth ( N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, 
        N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, 
        N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, 
        N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, 
        N74, N75, N76, N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, 
        N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, 
        N105, N106, N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, 
        N119, N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, 
        N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227, N230, 
        N231, N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, 
        N272, N275, N278, N281, N284, N287, N290, N294, N297, N301, N305, N309, 
        N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, 
        N349, N352, N355, N143_I, N144_I, N145_I, N146_I, N147_I, N148_I, 
        N149_I, N150_I, N151_I, N152_I, N153_I, N154_I, N155_I, N156_I, N157_I, 
        N158_I, N159_I, N160_I, N161_I, N162_I, N163_I, N164_I, N165_I, N166_I, 
        N167_I, N168_I, N169_I, N170_I, N171_I, N172_I, N173_I, N174_I, N175_I, 
        N176_I, N177_I, N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, 
        N185_I, N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I, 
        N194_I, N195_I, N196_I, N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, 
        N203_I, N204_I, N205_I, N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, 
        N212_I, N213_I, N214_I, N215_I, N216_I, N217_I, N218_I, N398, N400, 
        N401, N419, N420, N456, N457, N458, N487, N488, N489, N490, N491, N492, 
        N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, 
        N1726, N1816, N1817, N1818, N1819, N1820, N1821, N1969, N1970, N1971, 
        N2010, N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, 
        N2390, N2496, N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, 
        N3546, N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882, N143_O, 
        N144_O, N145_O, N146_O, N147_O, N148_O, N149_O, N150_O, N151_O, N152_O, 
        N153_O, N154_O, N155_O, N156_O, N157_O, N158_O, N159_O, N160_O, N161_O, 
        N162_O, N163_O, N164_O, N165_O, N166_O, N167_O, N168_O, N169_O, N170_O, 
        N171_O, N172_O, N173_O, N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, 
        N180_O, N181_O, N182_O, N183_O, N184_O, N185_O, N186_O, N187_O, N188_O, 
        N189_O, N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O, 
        N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O, N206_O, 
        N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, N214_O, N215_O, 
        N216_O, N217_O, N218_O );
  input N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40,
         N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119,
         N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227,
         N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263,
         N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297,
         N301, N305, N309, N313, N316, N319, N322, N325, N328, N331, N334,
         N337, N340, N343, N346, N349, N352, N355, N143_I, N144_I, N145_I,
         N146_I, N147_I, N148_I, N149_I, N150_I, N151_I, N152_I, N153_I,
         N154_I, N155_I, N156_I, N157_I, N158_I, N159_I, N160_I, N161_I,
         N162_I, N163_I, N164_I, N165_I, N166_I, N167_I, N168_I, N169_I,
         N170_I, N171_I, N172_I, N173_I, N174_I, N175_I, N176_I, N177_I,
         N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, N185_I,
         N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I,
         N194_I, N195_I, N196_I, N197_I, N198_I, N199_I, N200_I, N201_I,
         N202_I, N203_I, N204_I, N205_I, N206_I, N207_I, N208_I, N209_I,
         N210_I, N211_I, N212_I, N213_I, N214_I, N215_I, N216_I, N217_I,
         N218_I;
  output N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489,
         N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029,
         N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821,
         N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022,
         N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970,
         N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875,
         N3881, N3882, N143_O, N144_O, N145_O, N146_O, N147_O, N148_O, N149_O,
         N150_O, N151_O, N152_O, N153_O, N154_O, N155_O, N156_O, N157_O,
         N158_O, N159_O, N160_O, N161_O, N162_O, N163_O, N164_O, N165_O,
         N166_O, N167_O, N168_O, N169_O, N170_O, N171_O, N172_O, N173_O,
         N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, N180_O, N181_O,
         N182_O, N183_O, N184_O, N185_O, N186_O, N187_O, N188_O, N189_O,
         N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O,
         N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O,
         N206_O, N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, N213_O,
         N214_O, N215_O, N216_O, N217_O, N218_O;
  wire   N405, N408, N425, N485, N486, N495, N496, N499, N500, N503, N506,
         N509, N521, N533, N537, N543, N544, N547, N550, N562, N574, N578,
         N582, N594, N606, N607, N608, N609, N610, N611, N612, N613, N625,
         N637, N643, N650, N651, N655, N659, N663, N667, N671, N675, N679,
         N683, N687, N693, N699, N705, N711, N715, N719, N723, N727, N730,
         N733, N734, N735, N738, N741, N744, N747, N750, N753, N756, N759,
         N762, N765, N768, N771, N774, N777, N780, N783, N786, N800, N900,
         N901, N902, N903, N904, N905, N998, N999, N1027, N1032, N1033, N1034,
         N1037, N1042, N1053, N1064, N1065, N1066, N1067, N1068, N1069, N1070,
         N1075, N1086, N1097, N1098, N1099, N1100, N1101, N1102, N1113, N1124,
         N1125, N1126, N1127, N1128, N1129, N1133, N1137, N1140, N1141, N1142,
         N1143, N1144, N1145, N1146, N1157, N1168, N1169, N1170, N1171, N1172,
         N1173, N1178, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1195,
         N1200, N1205, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1219,
         N1222, N1225, N1228, N1231, N1234, N1237, N1240, N1243, N1246, N1249,
         N1250, N1251, N1254, N1257, N1260, N1263, N1266, N1275, N1276, N1302,
         N1351, N1352, N1353, N1354, N1355, N1395, N1396, N1397, N1398, N1399,
         N1422, N1423, N1424, N1425, N1426, N1427, N1440, N1441, N1449, N1450,
         N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460,
         N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470,
         N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480,
         N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490,
         N1491, N1492, N1493, N1494, N1495, N1496, N1499, N1502, N1506, N1510,
         N1513, N1516, N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526,
         N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536,
         N1537, N1538, N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546,
         N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1557, N1561, N1564,
         N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573, N1574,
         N1575, N1576, N1577, N1578, N1581, N1582, N1585, N1588, N1591, N1596,
         N1600, N1606, N1612, N1615, N1619, N1624, N1628, N1631, N1634, N1637,
         N1642, N1647, N1651, N1656, N1676, N1681, N1686, N1690, N1708, N1770,
         N1773, N1776, N1777, N1778, N1781, N1784, N1785, N1795, N1798, N1801,
         N1804, N1807, N1808, N1809, N1810, N1811, N1813, N1814, N1815, N1822,
         N1823, N1824, N1827, N1830, N1831, N1832, N1833, N1836, N1841, N1848,
         N1852, N1856, N1863, N1870, N1875, N1880, N1885, N1888, N1891, N1894,
         N1897, N1908, N1909, N1910, N1911, N1912, N1913, N1914, N1915, N1916,
         N1917, N1918, N1919, N1928, N1929, N1930, N1931, N1932, N1933, N1934,
         N1935, N1936, N1939, N1940, N1941, N1942, N1945, N1948, N1951, N1954,
         N1957, N1960, N1963, N1966, N2028, N2029, N2030, N2031, N2032, N2033,
         N2034, N2040, N2041, N2042, N2043, N2046, N2049, N2052, N2055, N2058,
         N2061, N2064, N2067, N2070, N2073, N2076, N2079, N2095, N2098, N2101,
         N2104, N2107, N2110, N2113, N2119, N2120, N2125, N2126, N2127, N2128,
         N2135, N2141, N2144, N2147, N2150, N2153, N2154, N2155, N2156, N2157,
         N2158, N2171, N2172, N2173, N2174, N2175, N2176, N2177, N2178, N2185,
         N2188, N2191, N2194, N2197, N2200, N2201, N2204, N2207, N2210, N2213,
         N2216, N2219, N2234, N2235, N2236, N2237, N2250, N2266, N2269, N2291,
         N2294, N2297, N2298, N2300, N2301, N2302, N2303, N2304, N2305, N2306,
         N2307, N2308, N2309, N2310, N2311, N2312, N2313, N2314, N2315, N2316,
         N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324, N2325, N2326,
         N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336,
         N2337, N2338, N2339, N2340, N2354, N2355, N2356, N2357, N2358, N2359,
         N2364, N2365, N2366, N2367, N2368, N2372, N2373, N2374, N2375, N2376,
         N2377, N2382, N2386, N2391, N2395, N2400, N2403, N2406, N2407, N2408,
         N2409, N2410, N2411, N2412, N2413, N2414, N2415, N2416, N2417, N2421,
         N2425, N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2437, N2440,
         N2443, N2446, N2449, N2452, N2453, N2454, N2457, N2460, N2463, N2466,
         N2469, N2472, N2475, N2478, N2481, N2484, N2487, N2490, N2493, N2503,
         N2504, N2510, N2511, N2521, N2528, N2531, N2534, N2537, N2540, N2544,
         N2545, N2546, N2547, N2548, N2549, N2550, N2551, N2552, N2553, N2563,
         N2564, N2565, N2566, N2567, N2568, N2579, N2603, N2607, N2608, N2609,
         N2610, N2611, N2612, N2613, N2617, N2618, N2619, N2620, N2621, N2624,
         N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2638,
         N2645, N2646, N2652, N2655, N2656, N2659, N2663, N2664, N2665, N2666,
         N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676,
         N2677, N2678, N2679, N2680, N2681, N2684, N2687, N2690, N2693, N2694,
         N2695, N2696, N2697, N2698, N2699, N2700, N2701, N2702, N2703, N2706,
         N2707, N2708, N2709, N2710, N2719, N2720, N2726, N2729, N2738, N2743,
         N2747, N2748, N2749, N2750, N2751, N2760, N2761, N2766, N2771, N2772,
         N2773, N2774, N2775, N2776, N2777, N2778, N2781, N2782, N2783, N2784,
         N2789, N2790, N2791, N2792, N2793, N2796, N2800, N2803, N2806, N2809,
         N2810, N2811, N2812, N2817, N2820, N2826, N2829, N2830, N2831, N2837,
         N2838, N2839, N2840, N2841, N2844, N2854, N2859, N2869, N2874, N2877,
         N2880, N2881, N2882, N2885, N2888, N2894, N2895, N2896, N2897, N2898,
         N2899, N2900, N2901, N2914, N2915, N2916, N2917, N2918, N2919, N2920,
         N2921, N2931, N2938, N2939, N2963, N2972, N2975, N2978, N2981, N2984,
         N2985, N2986, N2989, N2992, N2995, N2998, N3001, N3004, N3007, N3008,
         N3009, N3010, N3013, N3016, N3019, N3022, N3025, N3028, N3029, N3030,
         N3035, N3036, N3037, N3039, N3044, N3045, N3046, N3047, N3048, N3049,
         N3050, N3053, N3054, N3055, N3056, N3057, N3058, N3059, N3060, N3061,
         N3064, N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073,
         N3074, N3075, N3076, N3088, N3091, N3110, N3113, N3137, N3140, N3143,
         N3146, N3149, N3152, N3157, N3160, N3163, N3166, N3169, N3172, N3175,
         N3176, N3177, N3178, N3180, N3187, N3188, N3189, N3190, N3191, N3192,
         N3193, N3194, N3195, N3196, N3197, N3208, N3215, N3216, N3217, N3218,
         N3219, N3220, N3222, N3223, N3230, N3231, N3238, N3241, N3244, N3247,
         N3250, N3253, N3256, N3259, N3262, N3265, N3268, N3271, N3274, N3277,
         N3281, N3282, N3283, N3284, N3286, N3288, N3289, N3291, N3293, N3295,
         N3296, N3299, N3301, N3302, N3304, N3306, N3308, N3309, N3312, N3314,
         N3315, N3318, N3321, N3324, N3327, N3330, N3333, N3334, N3335, N3336,
         N3337, N3340, N3344, N3348, N3352, N3356, N3360, N3364, N3367, N3370,
         N3374, N3378, N3382, N3386, N3390, N3394, N3397, N3400, N3401, N3402,
         N3403, N3404, N3405, N3406, N3409, N3410, N3412, N3414, N3416, N3418,
         N3420, N3422, N3428, N3430, N3432, N3434, N3436, N3438, N3440, N3450,
         N3453, N3456, N3459, N3478, N3479, N3480, N3481, N3482, N3483, N3484,
         N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3494,
         N3496, N3498, N3499, N3500, N3501, N3502, N3503, N3504, N3505, N3506,
         N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3515, N3517, N3522,
         N3525, N3528, N3531, N3534, N3537, N3540, N3543, N3551, N3552, N3553,
         N3554, N3555, N3556, N3557, N3558, N3559, N3563, N3564, N3565, N3566,
         N3567, N3568, N3569, N3570, N3576, N3579, N3585, N3588, N3592, N3593,
         N3594, N3595, N3596, N3597, N3598, N3599, N3600, N3603, N3608, N3612,
         N3615, N3616, N3622, N3629, N3630, N3631, N3632, N3633, N3634, N3635,
         N3640, N3644, N3647, N3648, N3654, N3661, N3662, N3667, N3668, N3669,
         N3670, N3691, N3692, N3693, N3694, N3695, N3696, N3697, N3716, N3717,
         N3718, N3719, N3720, N3721, N3722, N3723, N3726, N3727, N3728, N3729,
         N3730, N3731, N3732, N3733, N3734, N3735, N3736, N3737, N3740, N3741,
         N3742, N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3753,
         N3754, N3758, N3761, N3762, N3767, N3771, N3774, N3775, N3778, N3779,
         N3780, N3790, N3793, N3794, N3802, N3805, N3806, N3807, N3808, N3811,
         N3812, N3813, N3814, N3815, N3816, N3817, N3818, N3819, N3820, N3821,
         N3822, N3823, N3826, N3827, N3834, N3835, N3836, N3837, N3838, N3839,
         N3840, N3843, N3852, N3857, N3858, N3859, N3864, N3869, N3870, N3876,
         N3877, N485_1, N485_2, N495_1, N544_1, N544_2, N547_1, N547_2,
         N1064_1, N1065_1, N1066_1, N1067_1, N1068_1, N1097_1, N1098_1,
         N1099_1, N1100_1, N1101_1, N1124_1, N1125_1, N1126_1, N1127_1,
         N1168_1, N1169_1, N1170_1, N1171_1, N1172_1, N1451_1, N1452_1,
         N1453_1, N1454_1, N1455_1, N1456_1, N1457_1, N1458_1, N1459_1,
         N1460_1, N1461_1, N1462_1, N1463_1, N1464_1, N1465_1, N1466_1,
         N1467_1, N1468_1, N1469_1, N1470_1, N1471_1, N1472_1, N1473_1,
         N1475_1, N1476_1, N1477_1, N1478_1, N1479_1, N1480_1, N1481_1,
         N1482_1, N1483_1, N1484_1, N1485_1, N1486_1, N1487_1, N1488_1,
         N1489_1, N1490_1, N1491_1, N1492_1, N1529_1, N1530_1, N1531_1,
         N1532_1, N1533_1, N1534_1, N1535_1, N1536_1, N1537_1, N1538_1,
         N1539_1, N1540_1, N1541_1, N1542_1, N1543_1, N1596_1, N1596_2,
         N1600_1, N1600_2, N1606_1, N1606_2, N1612_1, N1612_2, N1615_1,
         N1615_2, N1619_1, N1619_2, N1624_1, N1624_2, N1628_1, N1628_2,
         N1631_1, N1631_2, N1634_1, N1634_2, N1637_1, N1637_2, N1642_1,
         N1642_2, N1647_1, N1647_2, N1651_1, N1651_2, N1656_1, N1656_2,
         N1676_1, N1676_2, N1681_1, N1681_2, N1686_1, N1686_2, N1690_1,
         N1690_2, N1708_1, N1708_2, N1784_1, N1785_1, N1822_1, N1822_2,
         N1823_1, N1823_2, N1908_1, N1909_1, N2032_1, N2033_1, N2042_1,
         N2043_1, N2113_1, N2157_1, N2158_1, N2177_1, N2178_1, N2250_1,
         N2748_1, N2748_2, N2748_3, N2749_1, N2749_2, N2749_3, N2751_1,
         N2751_2, N2751_3, N2839_1, N2840_1, N2931_1, N2938_1, N2939_1,
         N3191_1, N3192_1, N3193_1, N3194_1, N3281_1, N3282_1, N3283_1,
         N3284_1, N3731_1, N3731_2, N3733_1, N3734_1, N3734_2, N3736_1,
         N3744_1, N3744_2, N3746_1, N3747_1, N3747_2, N3749_1, N3762_1,
         N3762_2, N3775_1, N3775_2, N3779_1, N3794_1, N3802_1, N3806_1,
         N3806_2, N3806_3, N3807_1, N3807_2, N3808_1, N3808_2, N3808_3,
         N3811_1, N3813_1, N3813_2, N3813_3, N3814_1, N3814_2, N3815_1,
         N3815_2, N3815_3, N3816_1, N3816_2, N3816_3, N3820_1, N3820_2,
         N3820_3, N3826_1, N3876_1, N3877_1;

  BUFX2 gate1 ( .A(N219), .Y(N398) );
  BUFX2 gate2 ( .A(N219), .Y(N400) );
  BUFX2 gate3 ( .A(N219), .Y(N401) );
  AND2X1 gate4 ( .A(N1), .B(N3), .Y(N405) );
  INVX1 gate5 ( .A(N230), .Y(N408) );
  BUFX2 gate6 ( .A(N253), .Y(N419) );
  BUFX2 gate7 ( .A(N253), .Y(N420) );
  INVX1 gate8 ( .A(N262), .Y(N425) );
  BUFX2 gate9 ( .A(N290), .Y(N456) );
  BUFX2 gate10 ( .A(N290), .Y(N457) );
  BUFX2 gate11 ( .A(N290), .Y(N458) );
  AND2X1 gate12_1 ( .A(N309), .B(N305), .Y(N485_1) );
  AND2X1 gate12_2 ( .A(N301), .B(N297), .Y(N485_2) );
  AND2X1 gate12 ( .A(N485_1), .B(N485_2), .Y(N485) );
  INVX1 gate13 ( .A(N405), .Y(N486) );
  INVX1 gate14 ( .A(N44), .Y(N487) );
  INVX1 gate15 ( .A(N132), .Y(N488) );
  INVX1 gate16 ( .A(N82), .Y(N489) );
  INVX1 gate17 ( .A(N96), .Y(N490) );
  INVX1 gate18 ( .A(N69), .Y(N491) );
  INVX1 gate19 ( .A(N120), .Y(N492) );
  INVX1 gate20 ( .A(N57), .Y(N493) );
  INVX1 gate21 ( .A(N108), .Y(N494) );
  AND2X1 gate22_1 ( .A(N2), .B(N15), .Y(N495_1) );
  AND2X1 gate22 ( .A(N237), .B(N495_1), .Y(N495) );
  BUFX2 gate23 ( .A(N237), .Y(N496) );
  AND2X1 gate24 ( .A(N37), .B(N37), .Y(N499) );
  BUFX2 gate25 ( .A(N219), .Y(N500) );
  BUFX2 gate26 ( .A(N8), .Y(N503) );
  BUFX2 gate27 ( .A(N8), .Y(N506) );
  BUFX2 gate28 ( .A(N227), .Y(N509) );
  BUFX2 gate29 ( .A(N234), .Y(N521) );
  INVX1 gate30 ( .A(N241), .Y(N533) );
  INVX1 gate31 ( .A(N246), .Y(N537) );
  AND2X1 gate32 ( .A(N11), .B(N246), .Y(N543) );
  AND2X1 gate33_1 ( .A(N132), .B(N82), .Y(N544_1) );
  AND2X1 gate33_2 ( .A(N96), .B(N44), .Y(N544_2) );
  AND2X1 gate33 ( .A(N544_1), .B(N544_2), .Y(N544) );
  AND2X1 gate34_1 ( .A(N120), .B(N57), .Y(N547_1) );
  AND2X1 gate34_2 ( .A(N108), .B(N69), .Y(N547_2) );
  AND2X1 gate34 ( .A(N547_1), .B(N547_2), .Y(N547) );
  BUFX2 gate35 ( .A(N227), .Y(N550) );
  BUFX2 gate36 ( .A(N234), .Y(N562) );
  INVX1 gate37 ( .A(N256), .Y(N574) );
  INVX1 gate38 ( .A(N259), .Y(N578) );
  BUFX2 gate39 ( .A(N319), .Y(N582) );
  BUFX2 gate40 ( .A(N322), .Y(N594) );
  INVX1 gate41 ( .A(N328), .Y(N606) );
  INVX1 gate42 ( .A(N331), .Y(N607) );
  INVX1 gate43 ( .A(N334), .Y(N608) );
  INVX1 gate44 ( .A(N337), .Y(N609) );
  INVX1 gate45 ( .A(N340), .Y(N610) );
  INVX1 gate46 ( .A(N343), .Y(N611) );
  INVX1 gate47 ( .A(N352), .Y(N612) );
  BUFX2 gate48 ( .A(N319), .Y(N613) );
  BUFX2 gate49 ( .A(N322), .Y(N625) );
  BUFX2 gate50 ( .A(N16), .Y(N637) );
  BUFX2 gate51 ( .A(N16), .Y(N643) );
  INVX1 gate52 ( .A(N355), .Y(N650) );
  AND2X1 gate53 ( .A(N7), .B(N237), .Y(N651) );
  INVX1 gate54 ( .A(N263), .Y(N655) );
  INVX1 gate55 ( .A(N266), .Y(N659) );
  INVX1 gate56 ( .A(N269), .Y(N663) );
  INVX1 gate57 ( .A(N272), .Y(N667) );
  INVX1 gate58 ( .A(N275), .Y(N671) );
  INVX1 gate59 ( .A(N278), .Y(N675) );
  INVX1 gate60 ( .A(N281), .Y(N679) );
  INVX1 gate61 ( .A(N284), .Y(N683) );
  INVX1 gate62 ( .A(N287), .Y(N687) );
  BUFX2 gate63 ( .A(N29), .Y(N693) );
  BUFX2 gate64 ( .A(N29), .Y(N699) );
  INVX1 gate65 ( .A(N294), .Y(N705) );
  INVX1 gate66 ( .A(N297), .Y(N711) );
  INVX1 gate67 ( .A(N301), .Y(N715) );
  INVX1 gate68 ( .A(N305), .Y(N719) );
  INVX1 gate69 ( .A(N309), .Y(N723) );
  INVX1 gate70 ( .A(N313), .Y(N727) );
  INVX1 gate71 ( .A(N316), .Y(N730) );
  INVX1 gate72 ( .A(N346), .Y(N733) );
  INVX1 gate73 ( .A(N349), .Y(N734) );
  BUFX2 gate74 ( .A(N259), .Y(N735) );
  BUFX2 gate75 ( .A(N256), .Y(N738) );
  BUFX2 gate76 ( .A(N263), .Y(N741) );
  BUFX2 gate77 ( .A(N269), .Y(N744) );
  BUFX2 gate78 ( .A(N266), .Y(N747) );
  BUFX2 gate79 ( .A(N275), .Y(N750) );
  BUFX2 gate80 ( .A(N272), .Y(N753) );
  BUFX2 gate81 ( .A(N281), .Y(N756) );
  BUFX2 gate82 ( .A(N278), .Y(N759) );
  BUFX2 gate83 ( .A(N287), .Y(N762) );
  BUFX2 gate84 ( .A(N284), .Y(N765) );
  BUFX2 gate85 ( .A(N294), .Y(N768) );
  BUFX2 gate86 ( .A(N301), .Y(N771) );
  BUFX2 gate87 ( .A(N297), .Y(N774) );
  BUFX2 gate88 ( .A(N309), .Y(N777) );
  BUFX2 gate89 ( .A(N305), .Y(N780) );
  BUFX2 gate90 ( .A(N316), .Y(N783) );
  BUFX2 gate91 ( .A(N313), .Y(N786) );
  INVX1 gate92 ( .A(N485), .Y(N792) );
  INVX1 gate93 ( .A(N495), .Y(N799) );
  INVX1 gate94 ( .A(N499), .Y(N800) );
  BUFX2 gate95 ( .A(N500), .Y(N805) );
  NAND2X1 gate96 ( .A(N331), .B(N606), .Y(N900) );
  NAND2X1 gate97 ( .A(N328), .B(N607), .Y(N901) );
  NAND2X1 gate98 ( .A(N337), .B(N608), .Y(N902) );
  NAND2X1 gate99 ( .A(N334), .B(N609), .Y(N903) );
  NAND2X1 gate100 ( .A(N343), .B(N610), .Y(N904) );
  NAND2X1 gate101 ( .A(N340), .B(N611), .Y(N905) );
  NAND2X1 gate102 ( .A(N349), .B(N733), .Y(N998) );
  NAND2X1 gate103 ( .A(N346), .B(N734), .Y(N999) );
  AND2X1 gate104 ( .A(N94), .B(N500), .Y(N1026) );
  AND2X1 gate105 ( .A(N325), .B(N651), .Y(N1027) );
  INVX1 gate106 ( .A(N651), .Y(N1028) );
  NAND2X1 gate107 ( .A(N231), .B(N651), .Y(N1029) );
  INVX1 gate108 ( .A(N544), .Y(N1032) );
  INVX1 gate109 ( .A(N547), .Y(N1033) );
  AND2X1 gate110 ( .A(N547), .B(N544), .Y(N1034) );
  BUFX2 gate111 ( .A(N503), .Y(N1037) );
  INVX1 gate112 ( .A(N509), .Y(N1042) );
  INVX1 gate113 ( .A(N521), .Y(N1053) );
  AND2X1 gate114_1 ( .A(N80), .B(N509), .Y(N1064_1) );
  AND2X1 gate114 ( .A(N521), .B(N1064_1), .Y(N1064) );
  AND2X1 gate115_1 ( .A(N68), .B(N509), .Y(N1065_1) );
  AND2X1 gate115 ( .A(N521), .B(N1065_1), .Y(N1065) );
  AND2X1 gate116_1 ( .A(N79), .B(N509), .Y(N1066_1) );
  AND2X1 gate116 ( .A(N521), .B(N1066_1), .Y(N1066) );
  AND2X1 gate117_1 ( .A(N78), .B(N509), .Y(N1067_1) );
  AND2X1 gate117 ( .A(N521), .B(N1067_1), .Y(N1067) );
  AND2X1 gate118_1 ( .A(N77), .B(N509), .Y(N1068_1) );
  AND2X1 gate118 ( .A(N521), .B(N1068_1), .Y(N1068) );
  AND2X1 gate119 ( .A(N11), .B(N537), .Y(N1069) );
  BUFX2 gate120 ( .A(N503), .Y(N1070) );
  INVX1 gate121 ( .A(N550), .Y(N1075) );
  INVX1 gate122 ( .A(N562), .Y(N1086) );
  AND2X1 gate123_1 ( .A(N76), .B(N550), .Y(N1097_1) );
  AND2X1 gate123 ( .A(N562), .B(N1097_1), .Y(N1097) );
  AND2X1 gate124_1 ( .A(N75), .B(N550), .Y(N1098_1) );
  AND2X1 gate124 ( .A(N562), .B(N1098_1), .Y(N1098) );
  AND2X1 gate125_1 ( .A(N74), .B(N550), .Y(N1099_1) );
  AND2X1 gate125 ( .A(N562), .B(N1099_1), .Y(N1099) );
  AND2X1 gate126_1 ( .A(N73), .B(N550), .Y(N1100_1) );
  AND2X1 gate126 ( .A(N562), .B(N1100_1), .Y(N1100) );
  AND2X1 gate127_1 ( .A(N72), .B(N550), .Y(N1101_1) );
  AND2X1 gate127 ( .A(N562), .B(N1101_1), .Y(N1101) );
  INVX1 gate128 ( .A(N582), .Y(N1102) );
  INVX1 gate129 ( .A(N594), .Y(N1113) );
  AND2X1 gate130_1 ( .A(N114), .B(N582), .Y(N1124_1) );
  AND2X1 gate130 ( .A(N594), .B(N1124_1), .Y(N1124) );
  AND2X1 gate131_1 ( .A(N113), .B(N582), .Y(N1125_1) );
  AND2X1 gate131 ( .A(N594), .B(N1125_1), .Y(N1125) );
  AND2X1 gate132_1 ( .A(N112), .B(N582), .Y(N1126_1) );
  AND2X1 gate132 ( .A(N594), .B(N1126_1), .Y(N1126) );
  AND2X1 gate133_1 ( .A(N111), .B(N582), .Y(N1127_1) );
  AND2X1 gate133 ( .A(N594), .B(N1127_1), .Y(N1127) );
  AND2X1 gate134 ( .A(N582), .B(N594), .Y(N1128) );
  NAND2X1 gate135 ( .A(N900), .B(N901), .Y(N1129) );
  NAND2X1 gate136 ( .A(N902), .B(N903), .Y(N1133) );
  NAND2X1 gate137 ( .A(N904), .B(N905), .Y(N1137) );
  INVX1 gate138 ( .A(N741), .Y(N1140) );
  NAND2X1 gate139 ( .A(N741), .B(N612), .Y(N1141) );
  INVX1 gate140 ( .A(N744), .Y(N1142) );
  INVX1 gate141 ( .A(N747), .Y(N1143) );
  INVX1 gate142 ( .A(N750), .Y(N1144) );
  INVX1 gate143 ( .A(N753), .Y(N1145) );
  INVX1 gate144 ( .A(N613), .Y(N1146) );
  INVX1 gate145 ( .A(N625), .Y(N1157) );
  AND2X1 gate146_1 ( .A(N118), .B(N613), .Y(N1168_1) );
  AND2X1 gate146 ( .A(N625), .B(N1168_1), .Y(N1168) );
  AND2X1 gate147_1 ( .A(N107), .B(N613), .Y(N1169_1) );
  AND2X1 gate147 ( .A(N625), .B(N1169_1), .Y(N1169) );
  AND2X1 gate148_1 ( .A(N117), .B(N613), .Y(N1170_1) );
  AND2X1 gate148 ( .A(N625), .B(N1170_1), .Y(N1170) );
  AND2X1 gate149_1 ( .A(N116), .B(N613), .Y(N1171_1) );
  AND2X1 gate149 ( .A(N625), .B(N1171_1), .Y(N1171) );
  AND2X1 gate150_1 ( .A(N115), .B(N613), .Y(N1172_1) );
  AND2X1 gate150 ( .A(N625), .B(N1172_1), .Y(N1172) );
  INVX1 gate151 ( .A(N637), .Y(N1173) );
  INVX1 gate152 ( .A(N643), .Y(N1178) );
  INVX1 gate153 ( .A(N768), .Y(N1184) );
  NAND2X1 gate154 ( .A(N768), .B(N650), .Y(N1185) );
  INVX1 gate155 ( .A(N771), .Y(N1186) );
  INVX1 gate156 ( .A(N774), .Y(N1187) );
  INVX1 gate157 ( .A(N777), .Y(N1188) );
  INVX1 gate158 ( .A(N780), .Y(N1189) );
  BUFX2 gate159 ( .A(N506), .Y(N1190) );
  BUFX2 gate160 ( .A(N506), .Y(N1195) );
  INVX1 gate161 ( .A(N693), .Y(N1200) );
  INVX1 gate162 ( .A(N699), .Y(N1205) );
  INVX1 gate163 ( .A(N735), .Y(N1210) );
  INVX1 gate164 ( .A(N738), .Y(N1211) );
  INVX1 gate165 ( .A(N756), .Y(N1212) );
  INVX1 gate166 ( .A(N759), .Y(N1213) );
  INVX1 gate167 ( .A(N762), .Y(N1214) );
  INVX1 gate168 ( .A(N765), .Y(N1215) );
  NAND2X1 gate169 ( .A(N998), .B(N999), .Y(N1216) );
  BUFX2 gate170 ( .A(N574), .Y(N1219) );
  BUFX2 gate171 ( .A(N578), .Y(N1222) );
  BUFX2 gate172 ( .A(N655), .Y(N1225) );
  BUFX2 gate173 ( .A(N659), .Y(N1228) );
  BUFX2 gate174 ( .A(N663), .Y(N1231) );
  BUFX2 gate175 ( .A(N667), .Y(N1234) );
  BUFX2 gate176 ( .A(N671), .Y(N1237) );
  BUFX2 gate177 ( .A(N675), .Y(N1240) );
  BUFX2 gate178 ( .A(N679), .Y(N1243) );
  BUFX2 gate179 ( .A(N683), .Y(N1246) );
  INVX1 gate180 ( .A(N783), .Y(N1249) );
  INVX1 gate181 ( .A(N786), .Y(N1250) );
  BUFX2 gate182 ( .A(N687), .Y(N1251) );
  BUFX2 gate183 ( .A(N705), .Y(N1254) );
  BUFX2 gate184 ( .A(N711), .Y(N1257) );
  BUFX2 gate185 ( .A(N715), .Y(N1260) );
  BUFX2 gate186 ( .A(N719), .Y(N1263) );
  BUFX2 gate187 ( .A(N723), .Y(N1266) );
  INVX1 gate188 ( .A(N1027), .Y(N1269) );
  AND2X1 gate189 ( .A(N325), .B(N1032), .Y(N1275) );
  AND2X1 gate190 ( .A(N231), .B(N1033), .Y(N1276) );
  BUFX2 gate191 ( .A(N1034), .Y(N1277) );
  OR2X1 gate192 ( .A(N1069), .B(N543), .Y(N1302) );
  NAND2X1 gate193 ( .A(N352), .B(N1140), .Y(N1351) );
  NAND2X1 gate194 ( .A(N747), .B(N1142), .Y(N1352) );
  NAND2X1 gate195 ( .A(N744), .B(N1143), .Y(N1353) );
  NAND2X1 gate196 ( .A(N753), .B(N1144), .Y(N1354) );
  NAND2X1 gate197 ( .A(N750), .B(N1145), .Y(N1355) );
  NAND2X1 gate198 ( .A(N355), .B(N1184), .Y(N1395) );
  NAND2X1 gate199 ( .A(N774), .B(N1186), .Y(N1396) );
  NAND2X1 gate200 ( .A(N771), .B(N1187), .Y(N1397) );
  NAND2X1 gate201 ( .A(N780), .B(N1188), .Y(N1398) );
  NAND2X1 gate202 ( .A(N777), .B(N1189), .Y(N1399) );
  NAND2X1 gate203 ( .A(N738), .B(N1210), .Y(N1422) );
  NAND2X1 gate204 ( .A(N735), .B(N1211), .Y(N1423) );
  NAND2X1 gate205 ( .A(N759), .B(N1212), .Y(N1424) );
  NAND2X1 gate206 ( .A(N756), .B(N1213), .Y(N1425) );
  NAND2X1 gate207 ( .A(N765), .B(N1214), .Y(N1426) );
  NAND2X1 gate208 ( .A(N762), .B(N1215), .Y(N1427) );
  NAND2X1 gate209 ( .A(N786), .B(N1249), .Y(N1440) );
  NAND2X1 gate210 ( .A(N783), .B(N1250), .Y(N1441) );
  INVX1 gate211 ( .A(N1034), .Y(N1448) );
  INVX1 gate212 ( .A(N1275), .Y(N1449) );
  INVX1 gate213 ( .A(N1276), .Y(N1450) );
  AND2X1 gate214_1 ( .A(N93), .B(N1042), .Y(N1451_1) );
  AND2X1 gate214 ( .A(N1053), .B(N1451_1), .Y(N1451) );
  AND2X1 gate215_1 ( .A(N55), .B(N509), .Y(N1452_1) );
  AND2X1 gate215 ( .A(N1053), .B(N1452_1), .Y(N1452) );
  AND2X1 gate216_1 ( .A(N67), .B(N1042), .Y(N1453_1) );
  AND2X1 gate216 ( .A(N521), .B(N1453_1), .Y(N1453) );
  AND2X1 gate217_1 ( .A(N81), .B(N1042), .Y(N1454_1) );
  AND2X1 gate217 ( .A(N1053), .B(N1454_1), .Y(N1454) );
  AND2X1 gate218_1 ( .A(N43), .B(N509), .Y(N1455_1) );
  AND2X1 gate218 ( .A(N1053), .B(N1455_1), .Y(N1455) );
  AND2X1 gate219_1 ( .A(N56), .B(N1042), .Y(N1456_1) );
  AND2X1 gate219 ( .A(N521), .B(N1456_1), .Y(N1456) );
  AND2X1 gate220_1 ( .A(N92), .B(N1042), .Y(N1457_1) );
  AND2X1 gate220 ( .A(N1053), .B(N1457_1), .Y(N1457) );
  AND2X1 gate221_1 ( .A(N54), .B(N509), .Y(N1458_1) );
  AND2X1 gate221 ( .A(N1053), .B(N1458_1), .Y(N1458) );
  AND2X1 gate222_1 ( .A(N66), .B(N1042), .Y(N1459_1) );
  AND2X1 gate222 ( .A(N521), .B(N1459_1), .Y(N1459) );
  AND2X1 gate223_1 ( .A(N91), .B(N1042), .Y(N1460_1) );
  AND2X1 gate223 ( .A(N1053), .B(N1460_1), .Y(N1460) );
  AND2X1 gate224_1 ( .A(N53), .B(N509), .Y(N1461_1) );
  AND2X1 gate224 ( .A(N1053), .B(N1461_1), .Y(N1461) );
  AND2X1 gate225_1 ( .A(N65), .B(N1042), .Y(N1462_1) );
  AND2X1 gate225 ( .A(N521), .B(N1462_1), .Y(N1462) );
  AND2X1 gate226_1 ( .A(N90), .B(N1042), .Y(N1463_1) );
  AND2X1 gate226 ( .A(N1053), .B(N1463_1), .Y(N1463) );
  AND2X1 gate227_1 ( .A(N52), .B(N509), .Y(N1464_1) );
  AND2X1 gate227 ( .A(N1053), .B(N1464_1), .Y(N1464) );
  AND2X1 gate228_1 ( .A(N64), .B(N1042), .Y(N1465_1) );
  AND2X1 gate228 ( .A(N521), .B(N1465_1), .Y(N1465) );
  AND2X1 gate229_1 ( .A(N89), .B(N1075), .Y(N1466_1) );
  AND2X1 gate229 ( .A(N1086), .B(N1466_1), .Y(N1466) );
  AND2X1 gate230_1 ( .A(N51), .B(N550), .Y(N1467_1) );
  AND2X1 gate230 ( .A(N1086), .B(N1467_1), .Y(N1467) );
  AND2X1 gate231_1 ( .A(N63), .B(N1075), .Y(N1468_1) );
  AND2X1 gate231 ( .A(N562), .B(N1468_1), .Y(N1468) );
  AND2X1 gate232_1 ( .A(N88), .B(N1075), .Y(N1469_1) );
  AND2X1 gate232 ( .A(N1086), .B(N1469_1), .Y(N1469) );
  AND2X1 gate233_1 ( .A(N50), .B(N550), .Y(N1470_1) );
  AND2X1 gate233 ( .A(N1086), .B(N1470_1), .Y(N1470) );
  AND2X1 gate234_1 ( .A(N62), .B(N1075), .Y(N1471_1) );
  AND2X1 gate234 ( .A(N562), .B(N1471_1), .Y(N1471) );
  AND2X1 gate235_1 ( .A(N87), .B(N1075), .Y(N1472_1) );
  AND2X1 gate235 ( .A(N1086), .B(N1472_1), .Y(N1472) );
  AND2X1 gate236_1 ( .A(N49), .B(N550), .Y(N1473_1) );
  AND2X1 gate236 ( .A(N1086), .B(N1473_1), .Y(N1473) );
  AND2X1 gate237 ( .A(N1075), .B(N562), .Y(N1474) );
  AND2X1 gate238_1 ( .A(N86), .B(N1075), .Y(N1475_1) );
  AND2X1 gate238 ( .A(N1086), .B(N1475_1), .Y(N1475) );
  AND2X1 gate239_1 ( .A(N48), .B(N550), .Y(N1476_1) );
  AND2X1 gate239 ( .A(N1086), .B(N1476_1), .Y(N1476) );
  AND2X1 gate240_1 ( .A(N61), .B(N1075), .Y(N1477_1) );
  AND2X1 gate240 ( .A(N562), .B(N1477_1), .Y(N1477) );
  AND2X1 gate241_1 ( .A(N85), .B(N1075), .Y(N1478_1) );
  AND2X1 gate241 ( .A(N1086), .B(N1478_1), .Y(N1478) );
  AND2X1 gate242_1 ( .A(N47), .B(N550), .Y(N1479_1) );
  AND2X1 gate242 ( .A(N1086), .B(N1479_1), .Y(N1479) );
  AND2X1 gate243_1 ( .A(N60), .B(N1075), .Y(N1480_1) );
  AND2X1 gate243 ( .A(N562), .B(N1480_1), .Y(N1480) );
  AND2X1 gate244_1 ( .A(N138), .B(N1102), .Y(N1481_1) );
  AND2X1 gate244 ( .A(N1113), .B(N1481_1), .Y(N1481) );
  AND2X1 gate245_1 ( .A(N102), .B(N582), .Y(N1482_1) );
  AND2X1 gate245 ( .A(N1113), .B(N1482_1), .Y(N1482) );
  AND2X1 gate246_1 ( .A(N126), .B(N1102), .Y(N1483_1) );
  AND2X1 gate246 ( .A(N594), .B(N1483_1), .Y(N1483) );
  AND2X1 gate247_1 ( .A(N137), .B(N1102), .Y(N1484_1) );
  AND2X1 gate247 ( .A(N1113), .B(N1484_1), .Y(N1484) );
  AND2X1 gate248_1 ( .A(N101), .B(N582), .Y(N1485_1) );
  AND2X1 gate248 ( .A(N1113), .B(N1485_1), .Y(N1485) );
  AND2X1 gate249_1 ( .A(N125), .B(N1102), .Y(N1486_1) );
  AND2X1 gate249 ( .A(N594), .B(N1486_1), .Y(N1486) );
  AND2X1 gate250_1 ( .A(N136), .B(N1102), .Y(N1487_1) );
  AND2X1 gate250 ( .A(N1113), .B(N1487_1), .Y(N1487) );
  AND2X1 gate251_1 ( .A(N100), .B(N582), .Y(N1488_1) );
  AND2X1 gate251 ( .A(N1113), .B(N1488_1), .Y(N1488) );
  AND2X1 gate252_1 ( .A(N124), .B(N1102), .Y(N1489_1) );
  AND2X1 gate252 ( .A(N594), .B(N1489_1), .Y(N1489) );
  AND2X1 gate253_1 ( .A(N135), .B(N1102), .Y(N1490_1) );
  AND2X1 gate253 ( .A(N1113), .B(N1490_1), .Y(N1490) );
  AND2X1 gate254_1 ( .A(N99), .B(N582), .Y(N1491_1) );
  AND2X1 gate254 ( .A(N1113), .B(N1491_1), .Y(N1491) );
  AND2X1 gate255_1 ( .A(N123), .B(N1102), .Y(N1492_1) );
  AND2X1 gate255 ( .A(N594), .B(N1492_1), .Y(N1492) );
  AND2X1 gate256 ( .A(N1102), .B(N1113), .Y(N1493) );
  AND2X1 gate257 ( .A(N582), .B(N1113), .Y(N1494) );
  AND2X1 gate258 ( .A(N1102), .B(N594), .Y(N1495) );
  INVX1 gate259 ( .A(N1129), .Y(N1496) );
  INVX1 gate260 ( .A(N1133), .Y(N1499) );
  NAND2X1 gate261 ( .A(N1351), .B(N1141), .Y(N1502) );
  NAND2X1 gate262 ( .A(N1352), .B(N1353), .Y(N1506) );
  NAND2X1 gate263 ( .A(N1354), .B(N1355), .Y(N1510) );
  BUFX2 gate264 ( .A(N1137), .Y(N1513) );
  BUFX2 gate265 ( .A(N1137), .Y(N1516) );
  INVX1 gate266 ( .A(N1219), .Y(N1519) );
  INVX1 gate267 ( .A(N1222), .Y(N1520) );
  INVX1 gate268 ( .A(N1225), .Y(N1521) );
  INVX1 gate269 ( .A(N1228), .Y(N1522) );
  INVX1 gate270 ( .A(N1231), .Y(N1523) );
  INVX1 gate271 ( .A(N1234), .Y(N1524) );
  INVX1 gate272 ( .A(N1237), .Y(N1525) );
  INVX1 gate273 ( .A(N1240), .Y(N1526) );
  INVX1 gate274 ( .A(N1243), .Y(N1527) );
  INVX1 gate275 ( .A(N1246), .Y(N1528) );
  AND2X1 gate276_1 ( .A(N142), .B(N1146), .Y(N1529_1) );
  AND2X1 gate276 ( .A(N1157), .B(N1529_1), .Y(N1529) );
  AND2X1 gate277_1 ( .A(N106), .B(N613), .Y(N1530_1) );
  AND2X1 gate277 ( .A(N1157), .B(N1530_1), .Y(N1530) );
  AND2X1 gate278_1 ( .A(N130), .B(N1146), .Y(N1531_1) );
  AND2X1 gate278 ( .A(N625), .B(N1531_1), .Y(N1531) );
  AND2X1 gate279_1 ( .A(N131), .B(N1146), .Y(N1532_1) );
  AND2X1 gate279 ( .A(N1157), .B(N1532_1), .Y(N1532) );
  AND2X1 gate280_1 ( .A(N95), .B(N613), .Y(N1533_1) );
  AND2X1 gate280 ( .A(N1157), .B(N1533_1), .Y(N1533) );
  AND2X1 gate281_1 ( .A(N119), .B(N1146), .Y(N1534_1) );
  AND2X1 gate281 ( .A(N625), .B(N1534_1), .Y(N1534) );
  AND2X1 gate282_1 ( .A(N141), .B(N1146), .Y(N1535_1) );
  AND2X1 gate282 ( .A(N1157), .B(N1535_1), .Y(N1535) );
  AND2X1 gate283_1 ( .A(N105), .B(N613), .Y(N1536_1) );
  AND2X1 gate283 ( .A(N1157), .B(N1536_1), .Y(N1536) );
  AND2X1 gate284_1 ( .A(N129), .B(N1146), .Y(N1537_1) );
  AND2X1 gate284 ( .A(N625), .B(N1537_1), .Y(N1537) );
  AND2X1 gate285_1 ( .A(N140), .B(N1146), .Y(N1538_1) );
  AND2X1 gate285 ( .A(N1157), .B(N1538_1), .Y(N1538) );
  AND2X1 gate286_1 ( .A(N104), .B(N613), .Y(N1539_1) );
  AND2X1 gate286 ( .A(N1157), .B(N1539_1), .Y(N1539) );
  AND2X1 gate287_1 ( .A(N128), .B(N1146), .Y(N1540_1) );
  AND2X1 gate287 ( .A(N625), .B(N1540_1), .Y(N1540) );
  AND2X1 gate288_1 ( .A(N139), .B(N1146), .Y(N1541_1) );
  AND2X1 gate288 ( .A(N1157), .B(N1541_1), .Y(N1541) );
  AND2X1 gate289_1 ( .A(N103), .B(N613), .Y(N1542_1) );
  AND2X1 gate289 ( .A(N1157), .B(N1542_1), .Y(N1542) );
  AND2X1 gate290_1 ( .A(N127), .B(N1146), .Y(N1543_1) );
  AND2X1 gate290 ( .A(N625), .B(N1543_1), .Y(N1543) );
  AND2X1 gate291 ( .A(N19), .B(N1173), .Y(N1544) );
  AND2X1 gate292 ( .A(N4), .B(N1173), .Y(N1545) );
  AND2X1 gate293 ( .A(N20), .B(N1173), .Y(N1546) );
  AND2X1 gate294 ( .A(N5), .B(N1173), .Y(N1547) );
  AND2X1 gate295 ( .A(N21), .B(N1178), .Y(N1548) );
  AND2X1 gate296 ( .A(N22), .B(N1178), .Y(N1549) );
  AND2X1 gate297 ( .A(N23), .B(N1178), .Y(N1550) );
  AND2X1 gate298 ( .A(N6), .B(N1178), .Y(N1551) );
  AND2X1 gate299 ( .A(N24), .B(N1178), .Y(N1552) );
  NAND2X1 gate300 ( .A(N1395), .B(N1185), .Y(N1553) );
  NAND2X1 gate301 ( .A(N1396), .B(N1397), .Y(N1557) );
  NAND2X1 gate302 ( .A(N1398), .B(N1399), .Y(N1561) );
  AND2X1 gate303 ( .A(N25), .B(N1200), .Y(N1564) );
  AND2X1 gate304 ( .A(N32), .B(N1200), .Y(N1565) );
  AND2X1 gate305 ( .A(N26), .B(N1200), .Y(N1566) );
  AND2X1 gate306 ( .A(N33), .B(N1200), .Y(N1567) );
  AND2X1 gate307 ( .A(N27), .B(N1205), .Y(N1568) );
  AND2X1 gate308 ( .A(N34), .B(N1205), .Y(N1569) );
  AND2X1 gate309 ( .A(N35), .B(N1205), .Y(N1570) );
  AND2X1 gate310 ( .A(N28), .B(N1205), .Y(N1571) );
  INVX1 gate311 ( .A(N1251), .Y(N1572) );
  INVX1 gate312 ( .A(N1254), .Y(N1573) );
  INVX1 gate313 ( .A(N1257), .Y(N1574) );
  INVX1 gate314 ( .A(N1260), .Y(N1575) );
  INVX1 gate315 ( .A(N1263), .Y(N1576) );
  INVX1 gate316 ( .A(N1266), .Y(N1577) );
  NAND2X1 gate317 ( .A(N1422), .B(N1423), .Y(N1578) );
  INVX1 gate318 ( .A(N1216), .Y(N1581) );
  NAND2X1 gate319 ( .A(N1426), .B(N1427), .Y(N1582) );
  NAND2X1 gate320 ( .A(N1424), .B(N1425), .Y(N1585) );
  NAND2X1 gate321 ( .A(N1440), .B(N1441), .Y(N1588) );
  AND2X1 gate322 ( .A(N1449), .B(N1450), .Y(N1591) );
  OR2X1 gate323_1 ( .A(N1451), .B(N1452), .Y(N1596_1) );
  OR2X1 gate323_2 ( .A(N1453), .B(N1064), .Y(N1596_2) );
  OR2X1 gate323 ( .A(N1596_1), .B(N1596_2), .Y(N1596) );
  OR2X1 gate324_1 ( .A(N1454), .B(N1455), .Y(N1600_1) );
  OR2X1 gate324_2 ( .A(N1456), .B(N1065), .Y(N1600_2) );
  OR2X1 gate324 ( .A(N1600_1), .B(N1600_2), .Y(N1600) );
  OR2X1 gate325_1 ( .A(N1457), .B(N1458), .Y(N1606_1) );
  OR2X1 gate325_2 ( .A(N1459), .B(N1066), .Y(N1606_2) );
  OR2X1 gate325 ( .A(N1606_1), .B(N1606_2), .Y(N1606) );
  OR2X1 gate326_1 ( .A(N1460), .B(N1461), .Y(N1612_1) );
  OR2X1 gate326_2 ( .A(N1462), .B(N1067), .Y(N1612_2) );
  OR2X1 gate326 ( .A(N1612_1), .B(N1612_2), .Y(N1612) );
  OR2X1 gate327_1 ( .A(N1463), .B(N1464), .Y(N1615_1) );
  OR2X1 gate327_2 ( .A(N1465), .B(N1068), .Y(N1615_2) );
  OR2X1 gate327 ( .A(N1615_1), .B(N1615_2), .Y(N1615) );
  OR2X1 gate328_1 ( .A(N1466), .B(N1467), .Y(N1619_1) );
  OR2X1 gate328_2 ( .A(N1468), .B(N1097), .Y(N1619_2) );
  OR2X1 gate328 ( .A(N1619_1), .B(N1619_2), .Y(N1619) );
  OR2X1 gate329_1 ( .A(N1469), .B(N1470), .Y(N1624_1) );
  OR2X1 gate329_2 ( .A(N1471), .B(N1098), .Y(N1624_2) );
  OR2X1 gate329 ( .A(N1624_1), .B(N1624_2), .Y(N1624) );
  OR2X1 gate330_1 ( .A(N1472), .B(N1473), .Y(N1628_1) );
  OR2X1 gate330_2 ( .A(N1474), .B(N1099), .Y(N1628_2) );
  OR2X1 gate330 ( .A(N1628_1), .B(N1628_2), .Y(N1628) );
  OR2X1 gate331_1 ( .A(N1475), .B(N1476), .Y(N1631_1) );
  OR2X1 gate331_2 ( .A(N1477), .B(N1100), .Y(N1631_2) );
  OR2X1 gate331 ( .A(N1631_1), .B(N1631_2), .Y(N1631) );
  OR2X1 gate332_1 ( .A(N1478), .B(N1479), .Y(N1634_1) );
  OR2X1 gate332_2 ( .A(N1480), .B(N1101), .Y(N1634_2) );
  OR2X1 gate332 ( .A(N1634_1), .B(N1634_2), .Y(N1634) );
  OR2X1 gate333_1 ( .A(N1481), .B(N1482), .Y(N1637_1) );
  OR2X1 gate333_2 ( .A(N1483), .B(N1124), .Y(N1637_2) );
  OR2X1 gate333 ( .A(N1637_1), .B(N1637_2), .Y(N1637) );
  OR2X1 gate334_1 ( .A(N1484), .B(N1485), .Y(N1642_1) );
  OR2X1 gate334_2 ( .A(N1486), .B(N1125), .Y(N1642_2) );
  OR2X1 gate334 ( .A(N1642_1), .B(N1642_2), .Y(N1642) );
  OR2X1 gate335_1 ( .A(N1487), .B(N1488), .Y(N1647_1) );
  OR2X1 gate335_2 ( .A(N1489), .B(N1126), .Y(N1647_2) );
  OR2X1 gate335 ( .A(N1647_1), .B(N1647_2), .Y(N1647) );
  OR2X1 gate336_1 ( .A(N1490), .B(N1491), .Y(N1651_1) );
  OR2X1 gate336_2 ( .A(N1492), .B(N1127), .Y(N1651_2) );
  OR2X1 gate336 ( .A(N1651_1), .B(N1651_2), .Y(N1651) );
  OR2X1 gate337_1 ( .A(N1493), .B(N1494), .Y(N1656_1) );
  OR2X1 gate337_2 ( .A(N1495), .B(N1128), .Y(N1656_2) );
  OR2X1 gate337 ( .A(N1656_1), .B(N1656_2), .Y(N1656) );
  OR2X1 gate338_1 ( .A(N1532), .B(N1533), .Y(N1676_1) );
  OR2X1 gate338_2 ( .A(N1534), .B(N1169), .Y(N1676_2) );
  OR2X1 gate338 ( .A(N1676_1), .B(N1676_2), .Y(N1676) );
  OR2X1 gate339_1 ( .A(N1535), .B(N1536), .Y(N1681_1) );
  OR2X1 gate339_2 ( .A(N1537), .B(N1170), .Y(N1681_2) );
  OR2X1 gate339 ( .A(N1681_1), .B(N1681_2), .Y(N1681) );
  OR2X1 gate340_1 ( .A(N1538), .B(N1539), .Y(N1686_1) );
  OR2X1 gate340_2 ( .A(N1540), .B(N1171), .Y(N1686_2) );
  OR2X1 gate340 ( .A(N1686_1), .B(N1686_2), .Y(N1686) );
  OR2X1 gate341_1 ( .A(N1541), .B(N1542), .Y(N1690_1) );
  OR2X1 gate341_2 ( .A(N1543), .B(N1172), .Y(N1690_2) );
  OR2X1 gate341 ( .A(N1690_1), .B(N1690_2), .Y(N1690) );
  OR2X1 gate342_1 ( .A(N1529), .B(N1530), .Y(N1708_1) );
  OR2X1 gate342_2 ( .A(N1531), .B(N1168), .Y(N1708_2) );
  OR2X1 gate342 ( .A(N1708_1), .B(N1708_2), .Y(N1708) );
  BUFX2 gate343 ( .A(N1591), .Y(N1726) );
  INVX1 gate344 ( .A(N1502), .Y(N1770) );
  INVX1 gate345 ( .A(N1506), .Y(N1773) );
  INVX1 gate346 ( .A(N1513), .Y(N1776) );
  INVX1 gate347 ( .A(N1516), .Y(N1777) );
  BUFX2 gate348 ( .A(N1510), .Y(N1778) );
  BUFX2 gate349 ( .A(N1510), .Y(N1781) );
  AND2X1 gate350_1 ( .A(N1133), .B(N1129), .Y(N1784_1) );
  AND2X1 gate350 ( .A(N1513), .B(N1784_1), .Y(N1784) );
  AND2X1 gate351_1 ( .A(N1499), .B(N1496), .Y(N1785_1) );
  AND2X1 gate351 ( .A(N1516), .B(N1785_1), .Y(N1785) );
  INVX1 gate352 ( .A(N1553), .Y(N1795) );
  INVX1 gate353 ( .A(N1557), .Y(N1798) );
  BUFX2 gate354 ( .A(N1561), .Y(N1801) );
  BUFX2 gate355 ( .A(N1561), .Y(N1804) );
  INVX1 gate356 ( .A(N1588), .Y(N1807) );
  INVX1 gate357 ( .A(N1578), .Y(N1808) );
  NAND2X1 gate358 ( .A(N1578), .B(N1581), .Y(N1809) );
  INVX1 gate359 ( .A(N1582), .Y(N1810) );
  INVX1 gate360 ( .A(N1585), .Y(N1811) );
  AND2X1 gate361 ( .A(N1596), .B(N241), .Y(N1813) );
  AND2X1 gate362 ( .A(N1606), .B(N241), .Y(N1814) );
  AND2X1 gate363 ( .A(N1600), .B(N241), .Y(N1815) );
  INVX1 gate364 ( .A(N1642), .Y(N1816) );
  INVX1 gate365 ( .A(N1647), .Y(N1817) );
  INVX1 gate366 ( .A(N1637), .Y(N1818) );
  INVX1 gate367 ( .A(N1624), .Y(N1819) );
  INVX1 gate368 ( .A(N1619), .Y(N1820) );
  INVX1 gate369 ( .A(N1615), .Y(N1821) );
  AND2X1 gate370_1 ( .A(N496), .B(N224), .Y(N1822_1) );
  AND2X1 gate370_2 ( .A(N36), .B(N1591), .Y(N1822_2) );
  AND2X1 gate370 ( .A(N1822_1), .B(N1822_2), .Y(N1822) );
  AND2X1 gate371_1 ( .A(N496), .B(N224), .Y(N1823_1) );
  AND2X1 gate371_2 ( .A(N1591), .B(N486), .Y(N1823_2) );
  AND2X1 gate371 ( .A(N1823_1), .B(N1823_2), .Y(N1823) );
  BUFX2 gate372 ( .A(N1596), .Y(N1824) );
  INVX1 gate373 ( .A(N1606), .Y(N1827) );
  AND2X1 gate374 ( .A(N1600), .B(N537), .Y(N1830) );
  AND2X1 gate375 ( .A(N1606), .B(N537), .Y(N1831) );
  AND2X1 gate376 ( .A(N1619), .B(N246), .Y(N1832) );
  INVX1 gate377 ( .A(N1596), .Y(N1833) );
  INVX1 gate378 ( .A(N1600), .Y(N1836) );
  INVX1 gate379 ( .A(N1606), .Y(N1841) );
  BUFX2 gate380 ( .A(N1612), .Y(N1848) );
  BUFX2 gate381 ( .A(N1615), .Y(N1852) );
  BUFX2 gate382 ( .A(N1619), .Y(N1856) );
  BUFX2 gate383 ( .A(N1624), .Y(N1863) );
  BUFX2 gate384 ( .A(N1628), .Y(N1870) );
  BUFX2 gate385 ( .A(N1631), .Y(N1875) );
  BUFX2 gate386 ( .A(N1634), .Y(N1880) );
  NAND2X1 gate387 ( .A(N727), .B(N1651), .Y(N1885) );
  NAND2X1 gate388 ( .A(N730), .B(N1656), .Y(N1888) );
  BUFX2 gate389 ( .A(N1686), .Y(N1891) );
  AND2X1 gate390 ( .A(N1637), .B(N425), .Y(N1894) );
  INVX1 gate391 ( .A(N1642), .Y(N1897) );
  AND2X1 gate392_1 ( .A(N1496), .B(N1133), .Y(N1908_1) );
  AND2X1 gate392 ( .A(N1776), .B(N1908_1), .Y(N1908) );
  AND2X1 gate393_1 ( .A(N1129), .B(N1499), .Y(N1909_1) );
  AND2X1 gate393 ( .A(N1777), .B(N1909_1), .Y(N1909) );
  AND2X1 gate394 ( .A(N1600), .B(N637), .Y(N1910) );
  AND2X1 gate395 ( .A(N1606), .B(N637), .Y(N1911) );
  AND2X1 gate396 ( .A(N1612), .B(N637), .Y(N1912) );
  AND2X1 gate397 ( .A(N1615), .B(N637), .Y(N1913) );
  AND2X1 gate398 ( .A(N1619), .B(N643), .Y(N1914) );
  AND2X1 gate399 ( .A(N1624), .B(N643), .Y(N1915) );
  AND2X1 gate400 ( .A(N1628), .B(N643), .Y(N1916) );
  AND2X1 gate401 ( .A(N1631), .B(N643), .Y(N1917) );
  AND2X1 gate402 ( .A(N1634), .B(N643), .Y(N1918) );
  INVX1 gate403 ( .A(N1708), .Y(N1919) );
  AND2X1 gate404 ( .A(N1676), .B(N693), .Y(N1928) );
  AND2X1 gate405 ( .A(N1681), .B(N693), .Y(N1929) );
  AND2X1 gate406 ( .A(N1686), .B(N693), .Y(N1930) );
  AND2X1 gate407 ( .A(N1690), .B(N693), .Y(N1931) );
  AND2X1 gate408 ( .A(N1637), .B(N699), .Y(N1932) );
  AND2X1 gate409 ( .A(N1642), .B(N699), .Y(N1933) );
  AND2X1 gate410 ( .A(N1647), .B(N699), .Y(N1934) );
  AND2X1 gate411 ( .A(N1651), .B(N699), .Y(N1935) );
  BUFX2 gate412 ( .A(N1600), .Y(N1936) );
  NAND2X1 gate413 ( .A(N1216), .B(N1808), .Y(N1939) );
  NAND2X1 gate414 ( .A(N1585), .B(N1810), .Y(N1940) );
  NAND2X1 gate415 ( .A(N1582), .B(N1811), .Y(N1941) );
  BUFX2 gate416 ( .A(N1676), .Y(N1942) );
  BUFX2 gate417 ( .A(N1686), .Y(N1945) );
  BUFX2 gate418 ( .A(N1681), .Y(N1948) );
  BUFX2 gate419 ( .A(N1637), .Y(N1951) );
  BUFX2 gate420 ( .A(N1690), .Y(N1954) );
  BUFX2 gate421 ( .A(N1647), .Y(N1957) );
  BUFX2 gate422 ( .A(N1642), .Y(N1960) );
  BUFX2 gate423 ( .A(N1656), .Y(N1963) );
  BUFX2 gate424 ( .A(N1651), .Y(N1966) );
  OR2X1 gate425 ( .A(N533), .B(N1815), .Y(N1969) );
  INVX1 gate426 ( .A(N1822), .Y(N1970) );
  INVX1 gate427 ( .A(N1823), .Y(N1971) );
  BUFX2 gate428 ( .A(N1848), .Y(N2010) );
  BUFX2 gate429 ( .A(N1852), .Y(N2012) );
  BUFX2 gate430 ( .A(N1856), .Y(N2014) );
  BUFX2 gate431 ( .A(N1863), .Y(N2016) );
  BUFX2 gate432 ( .A(N1870), .Y(N2018) );
  BUFX2 gate433 ( .A(N1875), .Y(N2020) );
  BUFX2 gate434 ( .A(N1880), .Y(N2022) );
  INVX1 gate435 ( .A(N1778), .Y(N2028) );
  INVX1 gate436 ( .A(N1781), .Y(N2029) );
  NOR2X1 gate437 ( .A(N1908), .B(N1784), .Y(N2030) );
  NOR2X1 gate438 ( .A(N1909), .B(N1785), .Y(N2031) );
  AND2X1 gate439_1 ( .A(N1506), .B(N1502), .Y(N2032_1) );
  AND2X1 gate439 ( .A(N1778), .B(N2032_1), .Y(N2032) );
  AND2X1 gate440_1 ( .A(N1773), .B(N1770), .Y(N2033_1) );
  AND2X1 gate440 ( .A(N1781), .B(N2033_1), .Y(N2033) );
  OR2X1 gate441 ( .A(N1571), .B(N1935), .Y(N2034) );
  INVX1 gate442 ( .A(N1801), .Y(N2040) );
  INVX1 gate443 ( .A(N1804), .Y(N2041) );
  AND2X1 gate444_1 ( .A(N1557), .B(N1553), .Y(N2042_1) );
  AND2X1 gate444 ( .A(N1801), .B(N2042_1), .Y(N2042) );
  AND2X1 gate445_1 ( .A(N1798), .B(N1795), .Y(N2043_1) );
  AND2X1 gate445 ( .A(N1804), .B(N2043_1), .Y(N2043) );
  NAND2X1 gate446 ( .A(N1939), .B(N1809), .Y(N2046) );
  NAND2X1 gate447 ( .A(N1940), .B(N1941), .Y(N2049) );
  OR2X1 gate448 ( .A(N1544), .B(N1910), .Y(N2052) );
  OR2X1 gate449 ( .A(N1545), .B(N1911), .Y(N2055) );
  OR2X1 gate450 ( .A(N1546), .B(N1912), .Y(N2058) );
  OR2X1 gate451 ( .A(N1547), .B(N1913), .Y(N2061) );
  OR2X1 gate452 ( .A(N1548), .B(N1914), .Y(N2064) );
  OR2X1 gate453 ( .A(N1549), .B(N1915), .Y(N2067) );
  OR2X1 gate454 ( .A(N1550), .B(N1916), .Y(N2070) );
  OR2X1 gate455 ( .A(N1551), .B(N1917), .Y(N2073) );
  OR2X1 gate456 ( .A(N1552), .B(N1918), .Y(N2076) );
  OR2X1 gate457 ( .A(N1564), .B(N1928), .Y(N2079) );
  OR2X1 gate458 ( .A(N1565), .B(N1929), .Y(N2095) );
  OR2X1 gate459 ( .A(N1566), .B(N1930), .Y(N2098) );
  OR2X1 gate460 ( .A(N1567), .B(N1931), .Y(N2101) );
  OR2X1 gate461 ( .A(N1568), .B(N1932), .Y(N2104) );
  OR2X1 gate462 ( .A(N1569), .B(N1933), .Y(N2107) );
  OR2X1 gate463 ( .A(N1570), .B(N1934), .Y(N2110) );
  AND2X1 gate464_1 ( .A(N1897), .B(N1894), .Y(N2113_1) );
  AND2X1 gate464 ( .A(N40), .B(N2113_1), .Y(N2113) );
  INVX1 gate465 ( .A(N1894), .Y(N2119) );
  NAND2X1 gate466 ( .A(N408), .B(N1827), .Y(N2120) );
  AND2X1 gate467 ( .A(N1824), .B(N537), .Y(N2125) );
  AND2X1 gate468 ( .A(N1852), .B(N246), .Y(N2126) );
  AND2X1 gate469 ( .A(N1848), .B(N537), .Y(N2127) );
  INVX1 gate470 ( .A(N1848), .Y(N2128) );
  INVX1 gate471 ( .A(N1852), .Y(N2135) );
  INVX1 gate472 ( .A(N1863), .Y(N2141) );
  INVX1 gate473 ( .A(N1870), .Y(N2144) );
  INVX1 gate474 ( .A(N1875), .Y(N2147) );
  INVX1 gate475 ( .A(N1880), .Y(N2150) );
  AND2X1 gate476 ( .A(N727), .B(N1885), .Y(N2153) );
  AND2X1 gate477 ( .A(N1885), .B(N1651), .Y(N2154) );
  AND2X1 gate478 ( .A(N730), .B(N1888), .Y(N2155) );
  AND2X1 gate479 ( .A(N1888), .B(N1656), .Y(N2156) );
  AND2X1 gate480_1 ( .A(N1770), .B(N1506), .Y(N2157_1) );
  AND2X1 gate480 ( .A(N2028), .B(N2157_1), .Y(N2157) );
  AND2X1 gate481_1 ( .A(N1502), .B(N1773), .Y(N2158_1) );
  AND2X1 gate481 ( .A(N2029), .B(N2158_1), .Y(N2158) );
  INVX1 gate482 ( .A(N1942), .Y(N2171) );
  NAND2X1 gate483 ( .A(N1942), .B(N1919), .Y(N2172) );
  INVX1 gate484 ( .A(N1945), .Y(N2173) );
  INVX1 gate485 ( .A(N1948), .Y(N2174) );
  INVX1 gate486 ( .A(N1951), .Y(N2175) );
  INVX1 gate487 ( .A(N1954), .Y(N2176) );
  AND2X1 gate488_1 ( .A(N1795), .B(N1557), .Y(N2177_1) );
  AND2X1 gate488 ( .A(N2040), .B(N2177_1), .Y(N2177) );
  AND2X1 gate489_1 ( .A(N1553), .B(N1798), .Y(N2178_1) );
  AND2X1 gate489 ( .A(N2041), .B(N2178_1), .Y(N2178) );
  BUFX2 gate490 ( .A(N1836), .Y(N2185) );
  BUFX2 gate491 ( .A(N1833), .Y(N2188) );
  BUFX2 gate492 ( .A(N1841), .Y(N2191) );
  INVX1 gate493 ( .A(N1856), .Y(N2194) );
  INVX1 gate494 ( .A(N1827), .Y(N2197) );
  INVX1 gate495 ( .A(N1936), .Y(N2200) );
  BUFX2 gate496 ( .A(N1836), .Y(N2201) );
  BUFX2 gate497 ( .A(N1833), .Y(N2204) );
  BUFX2 gate498 ( .A(N1841), .Y(N2207) );
  BUFX2 gate499 ( .A(N1824), .Y(N2210) );
  BUFX2 gate500 ( .A(N1841), .Y(N2213) );
  BUFX2 gate501 ( .A(N1841), .Y(N2216) );
  NAND2X1 gate502 ( .A(N2031), .B(N2030), .Y(N2219) );
  INVX1 gate503 ( .A(N1957), .Y(N2234) );
  INVX1 gate504 ( .A(N1960), .Y(N2235) );
  INVX1 gate505 ( .A(N1963), .Y(N2236) );
  INVX1 gate506 ( .A(N1966), .Y(N2237) );
  AND2X1 gate507_1 ( .A(N40), .B(N1897), .Y(N2250_1) );
  AND2X1 gate507 ( .A(N2119), .B(N2250_1), .Y(N2250) );
  OR2X1 gate508 ( .A(N1831), .B(N2126), .Y(N2266) );
  OR2X1 gate509 ( .A(N2127), .B(N1832), .Y(N2269) );
  OR2X1 gate510 ( .A(N2153), .B(N2154), .Y(N2291) );
  OR2X1 gate511 ( .A(N2155), .B(N2156), .Y(N2294) );
  NOR2X1 gate512 ( .A(N2157), .B(N2032), .Y(N2297) );
  NOR2X1 gate513 ( .A(N2158), .B(N2033), .Y(N2298) );
  INVX1 gate514 ( .A(N2046), .Y(N2300) );
  INVX1 gate515 ( .A(N2049), .Y(N2301) );
  NAND2X1 gate516 ( .A(N2052), .B(N1519), .Y(N2302) );
  INVX1 gate517 ( .A(N2052), .Y(N2303) );
  NAND2X1 gate518 ( .A(N2055), .B(N1520), .Y(N2304) );
  INVX1 gate519 ( .A(N2055), .Y(N2305) );
  NAND2X1 gate520 ( .A(N2058), .B(N1521), .Y(N2306) );
  INVX1 gate521 ( .A(N2058), .Y(N2307) );
  NAND2X1 gate522 ( .A(N2061), .B(N1522), .Y(N2308) );
  INVX1 gate523 ( .A(N2061), .Y(N2309) );
  NAND2X1 gate524 ( .A(N2064), .B(N1523), .Y(N2310) );
  INVX1 gate525 ( .A(N2064), .Y(N2311) );
  NAND2X1 gate526 ( .A(N2067), .B(N1524), .Y(N2312) );
  INVX1 gate527 ( .A(N2067), .Y(N2313) );
  NAND2X1 gate528 ( .A(N2070), .B(N1525), .Y(N2314) );
  INVX1 gate529 ( .A(N2070), .Y(N2315) );
  NAND2X1 gate530 ( .A(N2073), .B(N1526), .Y(N2316) );
  INVX1 gate531 ( .A(N2073), .Y(N2317) );
  NAND2X1 gate532 ( .A(N2076), .B(N1527), .Y(N2318) );
  INVX1 gate533 ( .A(N2076), .Y(N2319) );
  NAND2X1 gate534 ( .A(N2079), .B(N1528), .Y(N2320) );
  INVX1 gate535 ( .A(N2079), .Y(N2321) );
  NAND2X1 gate536 ( .A(N1708), .B(N2171), .Y(N2322) );
  NAND2X1 gate537 ( .A(N1948), .B(N2173), .Y(N2323) );
  NAND2X1 gate538 ( .A(N1945), .B(N2174), .Y(N2324) );
  NAND2X1 gate539 ( .A(N1954), .B(N2175), .Y(N2325) );
  NAND2X1 gate540 ( .A(N1951), .B(N2176), .Y(N2326) );
  NOR2X1 gate541 ( .A(N2177), .B(N2042), .Y(N2327) );
  NOR2X1 gate542 ( .A(N2178), .B(N2043), .Y(N2328) );
  NAND2X1 gate543 ( .A(N2095), .B(N1572), .Y(N2329) );
  INVX1 gate544 ( .A(N2095), .Y(N2330) );
  NAND2X1 gate545 ( .A(N2098), .B(N1573), .Y(N2331) );
  INVX1 gate546 ( .A(N2098), .Y(N2332) );
  NAND2X1 gate547 ( .A(N2101), .B(N1574), .Y(N2333) );
  INVX1 gate548 ( .A(N2101), .Y(N2334) );
  NAND2X1 gate549 ( .A(N2104), .B(N1575), .Y(N2335) );
  INVX1 gate550 ( .A(N2104), .Y(N2336) );
  NAND2X1 gate551 ( .A(N2107), .B(N1576), .Y(N2337) );
  INVX1 gate552 ( .A(N2107), .Y(N2338) );
  NAND2X1 gate553 ( .A(N2110), .B(N1577), .Y(N2339) );
  INVX1 gate554 ( .A(N2110), .Y(N2340) );
  NAND2X1 gate555 ( .A(N1960), .B(N2234), .Y(N2354) );
  NAND2X1 gate556 ( .A(N1957), .B(N2235), .Y(N2355) );
  NAND2X1 gate557 ( .A(N1966), .B(N2236), .Y(N2356) );
  NAND2X1 gate558 ( .A(N1963), .B(N2237), .Y(N2357) );
  AND2X1 gate559 ( .A(N2120), .B(N533), .Y(N2358) );
  INVX1 gate560 ( .A(N2113), .Y(N2359) );
  INVX1 gate561 ( .A(N2185), .Y(N2364) );
  INVX1 gate562 ( .A(N2188), .Y(N2365) );
  INVX1 gate563 ( .A(N2191), .Y(N2366) );
  INVX1 gate564 ( .A(N2194), .Y(N2367) );
  BUFX2 gate565 ( .A(N2120), .Y(N2368) );
  INVX1 gate566 ( .A(N2201), .Y(N2372) );
  INVX1 gate567 ( .A(N2204), .Y(N2373) );
  INVX1 gate568 ( .A(N2207), .Y(N2374) );
  INVX1 gate569 ( .A(N2210), .Y(N2375) );
  INVX1 gate570 ( .A(N2213), .Y(N2376) );
  INVX1 gate571 ( .A(N2113), .Y(N2377) );
  BUFX2 gate572 ( .A(N2113), .Y(N2382) );
  AND2X1 gate573 ( .A(N2120), .B(N246), .Y(N2386) );
  BUFX2 gate574 ( .A(N2266), .Y(N2387) );
  BUFX2 gate575 ( .A(N2266), .Y(N2388) );
  BUFX2 gate576 ( .A(N2269), .Y(N2389) );
  BUFX2 gate577 ( .A(N2269), .Y(N2390) );
  BUFX2 gate578 ( .A(N2113), .Y(N2391) );
  INVX1 gate579 ( .A(N2113), .Y(N2395) );
  NAND2X1 gate580 ( .A(N2219), .B(N2300), .Y(N2400) );
  INVX1 gate581 ( .A(N2216), .Y(N2403) );
  INVX1 gate582 ( .A(N2219), .Y(N2406) );
  NAND2X1 gate583 ( .A(N1219), .B(N2303), .Y(N2407) );
  NAND2X1 gate584 ( .A(N1222), .B(N2305), .Y(N2408) );
  NAND2X1 gate585 ( .A(N1225), .B(N2307), .Y(N2409) );
  NAND2X1 gate586 ( .A(N1228), .B(N2309), .Y(N2410) );
  NAND2X1 gate587 ( .A(N1231), .B(N2311), .Y(N2411) );
  NAND2X1 gate588 ( .A(N1234), .B(N2313), .Y(N2412) );
  NAND2X1 gate589 ( .A(N1237), .B(N2315), .Y(N2413) );
  NAND2X1 gate590 ( .A(N1240), .B(N2317), .Y(N2414) );
  NAND2X1 gate591 ( .A(N1243), .B(N2319), .Y(N2415) );
  NAND2X1 gate592 ( .A(N1246), .B(N2321), .Y(N2416) );
  NAND2X1 gate593 ( .A(N2322), .B(N2172), .Y(N2417) );
  NAND2X1 gate594 ( .A(N2323), .B(N2324), .Y(N2421) );
  NAND2X1 gate595 ( .A(N2325), .B(N2326), .Y(N2425) );
  NAND2X1 gate596 ( .A(N1251), .B(N2330), .Y(N2428) );
  NAND2X1 gate597 ( .A(N1254), .B(N2332), .Y(N2429) );
  NAND2X1 gate598 ( .A(N1257), .B(N2334), .Y(N2430) );
  NAND2X1 gate599 ( .A(N1260), .B(N2336), .Y(N2431) );
  NAND2X1 gate600 ( .A(N1263), .B(N2338), .Y(N2432) );
  NAND2X1 gate601 ( .A(N1266), .B(N2340), .Y(N2433) );
  BUFX2 gate602 ( .A(N2128), .Y(N2434) );
  BUFX2 gate603 ( .A(N2135), .Y(N2437) );
  BUFX2 gate604 ( .A(N2144), .Y(N2440) );
  BUFX2 gate605 ( .A(N2141), .Y(N2443) );
  BUFX2 gate606 ( .A(N2150), .Y(N2446) );
  BUFX2 gate607 ( .A(N2147), .Y(N2449) );
  INVX1 gate608 ( .A(N2197), .Y(N2452) );
  NAND2X1 gate609 ( .A(N2197), .B(N2200), .Y(N2453) );
  BUFX2 gate610 ( .A(N2128), .Y(N2454) );
  BUFX2 gate611 ( .A(N2144), .Y(N2457) );
  BUFX2 gate612 ( .A(N2141), .Y(N2460) );
  BUFX2 gate613 ( .A(N2150), .Y(N2463) );
  BUFX2 gate614 ( .A(N2147), .Y(N2466) );
  INVX1 gate615 ( .A(N2120), .Y(N2469) );
  BUFX2 gate616 ( .A(N2128), .Y(N2472) );
  BUFX2 gate617 ( .A(N2135), .Y(N2475) );
  BUFX2 gate618 ( .A(N2128), .Y(N2478) );
  BUFX2 gate619 ( .A(N2135), .Y(N2481) );
  NAND2X1 gate620 ( .A(N2298), .B(N2297), .Y(N2484) );
  NAND2X1 gate621 ( .A(N2356), .B(N2357), .Y(N2487) );
  NAND2X1 gate622 ( .A(N2354), .B(N2355), .Y(N2490) );
  NAND2X1 gate623 ( .A(N2328), .B(N2327), .Y(N2493) );
  OR2X1 gate624 ( .A(N2358), .B(N1814), .Y(N2496) );
  NAND2X1 gate625 ( .A(N2188), .B(N2364), .Y(N2503) );
  NAND2X1 gate626 ( .A(N2185), .B(N2365), .Y(N2504) );
  NAND2X1 gate627 ( .A(N2204), .B(N2372), .Y(N2510) );
  NAND2X1 gate628 ( .A(N2201), .B(N2373), .Y(N2511) );
  OR2X1 gate629 ( .A(N1830), .B(N2386), .Y(N2521) );
  NAND2X1 gate630 ( .A(N2046), .B(N2406), .Y(N2528) );
  INVX1 gate631 ( .A(N2291), .Y(N2531) );
  INVX1 gate632 ( .A(N2294), .Y(N2534) );
  BUFX2 gate633 ( .A(N2250), .Y(N2537) );
  BUFX2 gate634 ( .A(N2250), .Y(N2540) );
  NAND2X1 gate635 ( .A(N2302), .B(N2407), .Y(N2544) );
  NAND2X1 gate636 ( .A(N2304), .B(N2408), .Y(N2545) );
  NAND2X1 gate637 ( .A(N2306), .B(N2409), .Y(N2546) );
  NAND2X1 gate638 ( .A(N2308), .B(N2410), .Y(N2547) );
  NAND2X1 gate639 ( .A(N2310), .B(N2411), .Y(N2548) );
  NAND2X1 gate640 ( .A(N2312), .B(N2412), .Y(N2549) );
  NAND2X1 gate641 ( .A(N2314), .B(N2413), .Y(N2550) );
  NAND2X1 gate642 ( .A(N2316), .B(N2414), .Y(N2551) );
  NAND2X1 gate643 ( .A(N2318), .B(N2415), .Y(N2552) );
  NAND2X1 gate644 ( .A(N2320), .B(N2416), .Y(N2553) );
  NAND2X1 gate645 ( .A(N2329), .B(N2428), .Y(N2563) );
  NAND2X1 gate646 ( .A(N2331), .B(N2429), .Y(N2564) );
  NAND2X1 gate647 ( .A(N2333), .B(N2430), .Y(N2565) );
  NAND2X1 gate648 ( .A(N2335), .B(N2431), .Y(N2566) );
  NAND2X1 gate649 ( .A(N2337), .B(N2432), .Y(N2567) );
  NAND2X1 gate650 ( .A(N2339), .B(N2433), .Y(N2568) );
  NAND2X1 gate651 ( .A(N1936), .B(N2452), .Y(N2579) );
  BUFX2 gate652 ( .A(N2359), .Y(N2603) );
  AND2X1 gate653 ( .A(N1880), .B(N2377), .Y(N2607) );
  AND2X1 gate654 ( .A(N1676), .B(N2377), .Y(N2608) );
  AND2X1 gate655 ( .A(N1681), .B(N2377), .Y(N2609) );
  AND2X1 gate656 ( .A(N1891), .B(N2377), .Y(N2610) );
  AND2X1 gate657 ( .A(N1856), .B(N2382), .Y(N2611) );
  AND2X1 gate658 ( .A(N1863), .B(N2382), .Y(N2612) );
  NAND2X1 gate659 ( .A(N2503), .B(N2504), .Y(N2613) );
  INVX1 gate660 ( .A(N2434), .Y(N2617) );
  NAND2X1 gate661 ( .A(N2434), .B(N2366), .Y(N2618) );
  NAND2X1 gate662 ( .A(N2437), .B(N2367), .Y(N2619) );
  INVX1 gate663 ( .A(N2437), .Y(N2620) );
  INVX1 gate664 ( .A(N2368), .Y(N2621) );
  NAND2X1 gate665 ( .A(N2510), .B(N2511), .Y(N2624) );
  INVX1 gate666 ( .A(N2454), .Y(N2628) );
  NAND2X1 gate667 ( .A(N2454), .B(N2374), .Y(N2629) );
  INVX1 gate668 ( .A(N2472), .Y(N2630) );
  AND2X1 gate669 ( .A(N1856), .B(N2391), .Y(N2631) );
  AND2X1 gate670 ( .A(N1863), .B(N2391), .Y(N2632) );
  AND2X1 gate671 ( .A(N1880), .B(N2395), .Y(N2633) );
  AND2X1 gate672 ( .A(N1676), .B(N2395), .Y(N2634) );
  AND2X1 gate673 ( .A(N1681), .B(N2395), .Y(N2635) );
  AND2X1 gate674 ( .A(N1891), .B(N2395), .Y(N2636) );
  INVX1 gate675 ( .A(N2382), .Y(N2638) );
  BUFX2 gate676 ( .A(N2521), .Y(N2643) );
  BUFX2 gate677 ( .A(N2521), .Y(N2644) );
  INVX1 gate678 ( .A(N2475), .Y(N2645) );
  INVX1 gate679 ( .A(N2391), .Y(N2646) );
  NAND2X1 gate680 ( .A(N2528), .B(N2400), .Y(N2652) );
  INVX1 gate681 ( .A(N2478), .Y(N2655) );
  INVX1 gate682 ( .A(N2481), .Y(N2656) );
  BUFX2 gate683 ( .A(N2359), .Y(N2659) );
  INVX1 gate684 ( .A(N2484), .Y(N2663) );
  NAND2X1 gate685 ( .A(N2484), .B(N2301), .Y(N2664) );
  INVX1 gate686 ( .A(N2553), .Y(N2665) );
  INVX1 gate687 ( .A(N2552), .Y(N2666) );
  INVX1 gate688 ( .A(N2551), .Y(N2667) );
  INVX1 gate689 ( .A(N2550), .Y(N2668) );
  INVX1 gate690 ( .A(N2549), .Y(N2669) );
  INVX1 gate691 ( .A(N2548), .Y(N2670) );
  INVX1 gate692 ( .A(N2547), .Y(N2671) );
  INVX1 gate693 ( .A(N2546), .Y(N2672) );
  INVX1 gate694 ( .A(N2545), .Y(N2673) );
  INVX1 gate695 ( .A(N2544), .Y(N2674) );
  INVX1 gate696 ( .A(N2568), .Y(N2675) );
  INVX1 gate697 ( .A(N2567), .Y(N2676) );
  INVX1 gate698 ( .A(N2566), .Y(N2677) );
  INVX1 gate699 ( .A(N2565), .Y(N2678) );
  INVX1 gate700 ( .A(N2564), .Y(N2679) );
  INVX1 gate701 ( .A(N2563), .Y(N2680) );
  INVX1 gate702 ( .A(N2417), .Y(N2681) );
  INVX1 gate703 ( .A(N2421), .Y(N2684) );
  BUFX2 gate704 ( .A(N2425), .Y(N2687) );
  BUFX2 gate705 ( .A(N2425), .Y(N2690) );
  INVX1 gate706 ( .A(N2493), .Y(N2693) );
  NAND2X1 gate707 ( .A(N2493), .B(N1807), .Y(N2694) );
  INVX1 gate708 ( .A(N2440), .Y(N2695) );
  INVX1 gate709 ( .A(N2443), .Y(N2696) );
  INVX1 gate710 ( .A(N2446), .Y(N2697) );
  INVX1 gate711 ( .A(N2449), .Y(N2698) );
  INVX1 gate712 ( .A(N2457), .Y(N2699) );
  INVX1 gate713 ( .A(N2460), .Y(N2700) );
  INVX1 gate714 ( .A(N2463), .Y(N2701) );
  INVX1 gate715 ( .A(N2466), .Y(N2702) );
  NAND2X1 gate716 ( .A(N2579), .B(N2453), .Y(N2703) );
  INVX1 gate717 ( .A(N2469), .Y(N2706) );
  INVX1 gate718 ( .A(N2487), .Y(N2707) );
  INVX1 gate719 ( .A(N2490), .Y(N2708) );
  AND2X1 gate720 ( .A(N2294), .B(N2534), .Y(N2709) );
  AND2X1 gate721 ( .A(N2291), .B(N2531), .Y(N2710) );
  NAND2X1 gate722 ( .A(N2191), .B(N2617), .Y(N2719) );
  NAND2X1 gate723 ( .A(N2194), .B(N2620), .Y(N2720) );
  NAND2X1 gate724 ( .A(N2207), .B(N2628), .Y(N2726) );
  BUFX2 gate725 ( .A(N2537), .Y(N2729) );
  BUFX2 gate726 ( .A(N2537), .Y(N2738) );
  INVX1 gate727 ( .A(N2652), .Y(N2743) );
  NAND2X1 gate728 ( .A(N2049), .B(N2663), .Y(N2747) );
  AND2X1 gate729_1 ( .A(N2665), .B(N2666), .Y(N2748_1) );
  AND2X1 gate729_2 ( .A(N2667), .B(N2668), .Y(N2748_2) );
  AND2X1 gate729_3 ( .A(N2669), .B(N2748_1), .Y(N2748_3) );
  AND2X1 gate729 ( .A(N2748_2), .B(N2748_3), .Y(N2748) );
  AND2X1 gate730_1 ( .A(N2670), .B(N2671), .Y(N2749_1) );
  AND2X1 gate730_2 ( .A(N2672), .B(N2673), .Y(N2749_2) );
  AND2X1 gate730_3 ( .A(N2674), .B(N2749_1), .Y(N2749_3) );
  AND2X1 gate730 ( .A(N2749_2), .B(N2749_3), .Y(N2749) );
  AND2X1 gate731 ( .A(N2034), .B(N2675), .Y(N2750) );
  AND2X1 gate732_1 ( .A(N2676), .B(N2677), .Y(N2751_1) );
  AND2X1 gate732_2 ( .A(N2678), .B(N2679), .Y(N2751_2) );
  AND2X1 gate732_3 ( .A(N2680), .B(N2751_1), .Y(N2751_3) );
  AND2X1 gate732 ( .A(N2751_2), .B(N2751_3), .Y(N2751) );
  NAND2X1 gate733 ( .A(N1588), .B(N2693), .Y(N2760) );
  BUFX2 gate734 ( .A(N2540), .Y(N2761) );
  BUFX2 gate735 ( .A(N2540), .Y(N2766) );
  NAND2X1 gate736 ( .A(N2443), .B(N2695), .Y(N2771) );
  NAND2X1 gate737 ( .A(N2440), .B(N2696), .Y(N2772) );
  NAND2X1 gate738 ( .A(N2449), .B(N2697), .Y(N2773) );
  NAND2X1 gate739 ( .A(N2446), .B(N2698), .Y(N2774) );
  NAND2X1 gate740 ( .A(N2460), .B(N2699), .Y(N2775) );
  NAND2X1 gate741 ( .A(N2457), .B(N2700), .Y(N2776) );
  NAND2X1 gate742 ( .A(N2466), .B(N2701), .Y(N2777) );
  NAND2X1 gate743 ( .A(N2463), .B(N2702), .Y(N2778) );
  NAND2X1 gate744 ( .A(N2490), .B(N2707), .Y(N2781) );
  NAND2X1 gate745 ( .A(N2487), .B(N2708), .Y(N2782) );
  OR2X1 gate746 ( .A(N2709), .B(N2534), .Y(N2783) );
  OR2X1 gate747 ( .A(N2710), .B(N2531), .Y(N2784) );
  AND2X1 gate748 ( .A(N1856), .B(N2638), .Y(N2789) );
  AND2X1 gate749 ( .A(N1863), .B(N2638), .Y(N2790) );
  AND2X1 gate750 ( .A(N1870), .B(N2638), .Y(N2791) );
  AND2X1 gate751 ( .A(N1875), .B(N2638), .Y(N2792) );
  INVX1 gate752 ( .A(N2613), .Y(N2793) );
  NAND2X1 gate753 ( .A(N2719), .B(N2618), .Y(N2796) );
  NAND2X1 gate754 ( .A(N2619), .B(N2720), .Y(N2800) );
  INVX1 gate755 ( .A(N2624), .Y(N2803) );
  NAND2X1 gate756 ( .A(N2726), .B(N2629), .Y(N2806) );
  AND2X1 gate757 ( .A(N1856), .B(N2646), .Y(N2809) );
  AND2X1 gate758 ( .A(N1863), .B(N2646), .Y(N2810) );
  AND2X1 gate759 ( .A(N1870), .B(N2646), .Y(N2811) );
  AND2X1 gate760 ( .A(N1875), .B(N2646), .Y(N2812) );
  AND2X1 gate761 ( .A(N2743), .B(N14), .Y(N2817) );
  BUFX2 gate762 ( .A(N2603), .Y(N2820) );
  NAND2X1 gate763 ( .A(N2747), .B(N2664), .Y(N2826) );
  AND2X1 gate764 ( .A(N2748), .B(N2749), .Y(N2829) );
  AND2X1 gate765 ( .A(N2750), .B(N2751), .Y(N2830) );
  BUFX2 gate766 ( .A(N2659), .Y(N2831) );
  INVX1 gate767 ( .A(N2687), .Y(N2837) );
  INVX1 gate768 ( .A(N2690), .Y(N2838) );
  AND2X1 gate769_1 ( .A(N2421), .B(N2417), .Y(N2839_1) );
  AND2X1 gate769 ( .A(N2687), .B(N2839_1), .Y(N2839) );
  AND2X1 gate770_1 ( .A(N2684), .B(N2681), .Y(N2840_1) );
  AND2X1 gate770 ( .A(N2690), .B(N2840_1), .Y(N2840) );
  NAND2X1 gate771 ( .A(N2760), .B(N2694), .Y(N2841) );
  BUFX2 gate772 ( .A(N2603), .Y(N2844) );
  BUFX2 gate773 ( .A(N2603), .Y(N2854) );
  BUFX2 gate774 ( .A(N2659), .Y(N2859) );
  BUFX2 gate775 ( .A(N2659), .Y(N2869) );
  NAND2X1 gate776 ( .A(N2773), .B(N2774), .Y(N2874) );
  NAND2X1 gate777 ( .A(N2771), .B(N2772), .Y(N2877) );
  INVX1 gate778 ( .A(N2703), .Y(N2880) );
  NAND2X1 gate779 ( .A(N2703), .B(N2706), .Y(N2881) );
  NAND2X1 gate780 ( .A(N2777), .B(N2778), .Y(N2882) );
  NAND2X1 gate781 ( .A(N2775), .B(N2776), .Y(N2885) );
  NAND2X1 gate782 ( .A(N2781), .B(N2782), .Y(N2888) );
  NAND2X1 gate783 ( .A(N2783), .B(N2784), .Y(N2891) );
  AND2X1 gate784 ( .A(N2607), .B(N2729), .Y(N2894) );
  AND2X1 gate785 ( .A(N2608), .B(N2729), .Y(N2895) );
  AND2X1 gate786 ( .A(N2609), .B(N2729), .Y(N2896) );
  AND2X1 gate787 ( .A(N2610), .B(N2729), .Y(N2897) );
  OR2X1 gate788 ( .A(N2789), .B(N2611), .Y(N2898) );
  OR2X1 gate789 ( .A(N2790), .B(N2612), .Y(N2899) );
  AND2X1 gate790 ( .A(N2791), .B(N1037), .Y(N2900) );
  AND2X1 gate791 ( .A(N2792), .B(N1037), .Y(N2901) );
  OR2X1 gate792 ( .A(N2809), .B(N2631), .Y(N2914) );
  OR2X1 gate793 ( .A(N2810), .B(N2632), .Y(N2915) );
  AND2X1 gate794 ( .A(N2811), .B(N1070), .Y(N2916) );
  AND2X1 gate795 ( .A(N2812), .B(N1070), .Y(N2917) );
  AND2X1 gate796 ( .A(N2633), .B(N2738), .Y(N2918) );
  AND2X1 gate797 ( .A(N2634), .B(N2738), .Y(N2919) );
  AND2X1 gate798 ( .A(N2635), .B(N2738), .Y(N2920) );
  AND2X1 gate799 ( .A(N2636), .B(N2738), .Y(N2921) );
  BUFX2 gate800 ( .A(N2817), .Y(N2925) );
  AND2X1 gate801_1 ( .A(N2829), .B(N2830), .Y(N2931_1) );
  AND2X1 gate801 ( .A(N1302), .B(N2931_1), .Y(N2931) );
  AND2X1 gate802_1 ( .A(N2681), .B(N2421), .Y(N2938_1) );
  AND2X1 gate802 ( .A(N2837), .B(N2938_1), .Y(N2938) );
  AND2X1 gate803_1 ( .A(N2417), .B(N2684), .Y(N2939_1) );
  AND2X1 gate803 ( .A(N2838), .B(N2939_1), .Y(N2939) );
  NAND2X1 gate804 ( .A(N2469), .B(N2880), .Y(N2963) );
  INVX1 gate805 ( .A(N2841), .Y(N2970) );
  INVX1 gate806 ( .A(N2826), .Y(N2971) );
  INVX1 gate807 ( .A(N2894), .Y(N2972) );
  INVX1 gate808 ( .A(N2895), .Y(N2975) );
  INVX1 gate809 ( .A(N2896), .Y(N2978) );
  INVX1 gate810 ( .A(N2897), .Y(N2981) );
  AND2X1 gate811 ( .A(N2898), .B(N1037), .Y(N2984) );
  AND2X1 gate812 ( .A(N2899), .B(N1037), .Y(N2985) );
  INVX1 gate813 ( .A(N2900), .Y(N2986) );
  INVX1 gate814 ( .A(N2901), .Y(N2989) );
  INVX1 gate815 ( .A(N2796), .Y(N2992) );
  BUFX2 gate816 ( .A(N2800), .Y(N2995) );
  BUFX2 gate817 ( .A(N2800), .Y(N2998) );
  BUFX2 gate818 ( .A(N2806), .Y(N3001) );
  BUFX2 gate819 ( .A(N2806), .Y(N3004) );
  AND2X1 gate820 ( .A(N574), .B(N2820), .Y(N3007) );
  AND2X1 gate821 ( .A(N2914), .B(N1070), .Y(N3008) );
  AND2X1 gate822 ( .A(N2915), .B(N1070), .Y(N3009) );
  INVX1 gate823 ( .A(N2916), .Y(N3010) );
  INVX1 gate824 ( .A(N2917), .Y(N3013) );
  INVX1 gate825 ( .A(N2918), .Y(N3016) );
  INVX1 gate826 ( .A(N2919), .Y(N3019) );
  INVX1 gate827 ( .A(N2920), .Y(N3022) );
  INVX1 gate828 ( .A(N2921), .Y(N3025) );
  INVX1 gate829 ( .A(N2817), .Y(N3028) );
  AND2X1 gate830 ( .A(N574), .B(N2831), .Y(N3029) );
  INVX1 gate831 ( .A(N2820), .Y(N3030) );
  AND2X1 gate832 ( .A(N578), .B(N2820), .Y(N3035) );
  AND2X1 gate833 ( .A(N655), .B(N2820), .Y(N3036) );
  AND2X1 gate834 ( .A(N659), .B(N2820), .Y(N3037) );
  BUFX2 gate835 ( .A(N2931), .Y(N3038) );
  INVX1 gate836 ( .A(N2831), .Y(N3039) );
  AND2X1 gate837 ( .A(N578), .B(N2831), .Y(N3044) );
  AND2X1 gate838 ( .A(N655), .B(N2831), .Y(N3045) );
  AND2X1 gate839 ( .A(N659), .B(N2831), .Y(N3046) );
  NOR2X1 gate840 ( .A(N2938), .B(N2839), .Y(N3047) );
  NOR2X1 gate841 ( .A(N2939), .B(N2840), .Y(N3048) );
  INVX1 gate842 ( .A(N2888), .Y(N3049) );
  INVX1 gate843 ( .A(N2844), .Y(N3050) );
  AND2X1 gate844 ( .A(N663), .B(N2844), .Y(N3053) );
  AND2X1 gate845 ( .A(N667), .B(N2844), .Y(N3054) );
  AND2X1 gate846 ( .A(N671), .B(N2844), .Y(N3055) );
  AND2X1 gate847 ( .A(N675), .B(N2844), .Y(N3056) );
  AND2X1 gate848 ( .A(N679), .B(N2854), .Y(N3057) );
  AND2X1 gate849 ( .A(N683), .B(N2854), .Y(N3058) );
  AND2X1 gate850 ( .A(N687), .B(N2854), .Y(N3059) );
  AND2X1 gate851 ( .A(N705), .B(N2854), .Y(N3060) );
  INVX1 gate852 ( .A(N2859), .Y(N3061) );
  AND2X1 gate853 ( .A(N663), .B(N2859), .Y(N3064) );
  AND2X1 gate854 ( .A(N667), .B(N2859), .Y(N3065) );
  AND2X1 gate855 ( .A(N671), .B(N2859), .Y(N3066) );
  AND2X1 gate856 ( .A(N675), .B(N2859), .Y(N3067) );
  AND2X1 gate857 ( .A(N679), .B(N2869), .Y(N3068) );
  AND2X1 gate858 ( .A(N683), .B(N2869), .Y(N3069) );
  AND2X1 gate859 ( .A(N687), .B(N2869), .Y(N3070) );
  AND2X1 gate860 ( .A(N705), .B(N2869), .Y(N3071) );
  INVX1 gate861 ( .A(N2874), .Y(N3072) );
  INVX1 gate862 ( .A(N2877), .Y(N3073) );
  INVX1 gate863 ( .A(N2882), .Y(N3074) );
  INVX1 gate864 ( .A(N2885), .Y(N3075) );
  NAND2X1 gate865 ( .A(N2881), .B(N2963), .Y(N3076) );
  INVX1 gate866 ( .A(N2931), .Y(N3079) );
  INVX1 gate867 ( .A(N2984), .Y(N3088) );
  INVX1 gate868 ( .A(N2985), .Y(N3091) );
  INVX1 gate869 ( .A(N3008), .Y(N3110) );
  INVX1 gate870 ( .A(N3009), .Y(N3113) );
  AND2X1 gate871 ( .A(N3055), .B(N1190), .Y(N3137) );
  AND2X1 gate872 ( .A(N3056), .B(N1190), .Y(N3140) );
  AND2X1 gate873 ( .A(N3057), .B(N2761), .Y(N3143) );
  AND2X1 gate874 ( .A(N3058), .B(N2761), .Y(N3146) );
  AND2X1 gate875 ( .A(N3059), .B(N2761), .Y(N3149) );
  AND2X1 gate876 ( .A(N3060), .B(N2761), .Y(N3152) );
  AND2X1 gate877 ( .A(N3066), .B(N1195), .Y(N3157) );
  AND2X1 gate878 ( .A(N3067), .B(N1195), .Y(N3160) );
  AND2X1 gate879 ( .A(N3068), .B(N2766), .Y(N3163) );
  AND2X1 gate880 ( .A(N3069), .B(N2766), .Y(N3166) );
  AND2X1 gate881 ( .A(N3070), .B(N2766), .Y(N3169) );
  AND2X1 gate882 ( .A(N3071), .B(N2766), .Y(N3172) );
  NAND2X1 gate883 ( .A(N2877), .B(N3072), .Y(N3175) );
  NAND2X1 gate884 ( .A(N2874), .B(N3073), .Y(N3176) );
  NAND2X1 gate885 ( .A(N2885), .B(N3074), .Y(N3177) );
  NAND2X1 gate886 ( .A(N2882), .B(N3075), .Y(N3178) );
  NAND2X1 gate887 ( .A(N3048), .B(N3047), .Y(N3180) );
  INVX1 gate888 ( .A(N2995), .Y(N3187) );
  INVX1 gate889 ( .A(N2998), .Y(N3188) );
  INVX1 gate890 ( .A(N3001), .Y(N3189) );
  INVX1 gate891 ( .A(N3004), .Y(N3190) );
  AND2X1 gate892_1 ( .A(N2796), .B(N2613), .Y(N3191_1) );
  AND2X1 gate892 ( .A(N2995), .B(N3191_1), .Y(N3191) );
  AND2X1 gate893_1 ( .A(N2992), .B(N2793), .Y(N3192_1) );
  AND2X1 gate893 ( .A(N2998), .B(N3192_1), .Y(N3192) );
  AND2X1 gate894_1 ( .A(N2624), .B(N2368), .Y(N3193_1) );
  AND2X1 gate894 ( .A(N3001), .B(N3193_1), .Y(N3193) );
  AND2X1 gate895_1 ( .A(N2803), .B(N2621), .Y(N3194_1) );
  AND2X1 gate895 ( .A(N3004), .B(N3194_1), .Y(N3194) );
  NAND2X1 gate896 ( .A(N3076), .B(N2375), .Y(N3195) );
  INVX1 gate897 ( .A(N3076), .Y(N3196) );
  AND2X1 gate898 ( .A(N687), .B(N3030), .Y(N3197) );
  AND2X1 gate899 ( .A(N687), .B(N3039), .Y(N3208) );
  AND2X1 gate900 ( .A(N705), .B(N3030), .Y(N3215) );
  AND2X1 gate901 ( .A(N711), .B(N3030), .Y(N3216) );
  AND2X1 gate902 ( .A(N715), .B(N3030), .Y(N3217) );
  AND2X1 gate903 ( .A(N705), .B(N3039), .Y(N3218) );
  AND2X1 gate904 ( .A(N711), .B(N3039), .Y(N3219) );
  AND2X1 gate905 ( .A(N715), .B(N3039), .Y(N3220) );
  AND2X1 gate906 ( .A(N719), .B(N3050), .Y(N3222) );
  AND2X1 gate907 ( .A(N723), .B(N3050), .Y(N3223) );
  AND2X1 gate908 ( .A(N719), .B(N3061), .Y(N3230) );
  AND2X1 gate909 ( .A(N723), .B(N3061), .Y(N3231) );
  NAND2X1 gate910 ( .A(N3175), .B(N3176), .Y(N3238) );
  NAND2X1 gate911 ( .A(N3177), .B(N3178), .Y(N3241) );
  BUFX2 gate912 ( .A(N2981), .Y(N3244) );
  BUFX2 gate913 ( .A(N2978), .Y(N3247) );
  BUFX2 gate914 ( .A(N2975), .Y(N3250) );
  BUFX2 gate915 ( .A(N2972), .Y(N3253) );
  BUFX2 gate916 ( .A(N2989), .Y(N3256) );
  BUFX2 gate917 ( .A(N2986), .Y(N3259) );
  BUFX2 gate918 ( .A(N3025), .Y(N3262) );
  BUFX2 gate919 ( .A(N3022), .Y(N3265) );
  BUFX2 gate920 ( .A(N3019), .Y(N3268) );
  BUFX2 gate921 ( .A(N3016), .Y(N3271) );
  BUFX2 gate922 ( .A(N3013), .Y(N3274) );
  BUFX2 gate923 ( .A(N3010), .Y(N3277) );
  AND2X1 gate924_1 ( .A(N2793), .B(N2796), .Y(N3281_1) );
  AND2X1 gate924 ( .A(N3187), .B(N3281_1), .Y(N3281) );
  AND2X1 gate925_1 ( .A(N2613), .B(N2992), .Y(N3282_1) );
  AND2X1 gate925 ( .A(N3188), .B(N3282_1), .Y(N3282) );
  AND2X1 gate926_1 ( .A(N2621), .B(N2624), .Y(N3283_1) );
  AND2X1 gate926 ( .A(N3189), .B(N3283_1), .Y(N3283) );
  AND2X1 gate927_1 ( .A(N2368), .B(N2803), .Y(N3284_1) );
  AND2X1 gate927 ( .A(N3190), .B(N3284_1), .Y(N3284) );
  NAND2X1 gate928 ( .A(N2210), .B(N3196), .Y(N3286) );
  OR2X1 gate929 ( .A(N3197), .B(N3007), .Y(N3288) );
  NAND2X1 gate930 ( .A(N3180), .B(N3049), .Y(N3289) );
  AND2X1 gate931 ( .A(N3152), .B(N2981), .Y(N3291) );
  AND2X1 gate932 ( .A(N3149), .B(N2978), .Y(N3293) );
  AND2X1 gate933 ( .A(N3146), .B(N2975), .Y(N3295) );
  AND2X1 gate934 ( .A(N2972), .B(N3143), .Y(N3296) );
  AND2X1 gate935 ( .A(N3140), .B(N2989), .Y(N3299) );
  AND2X1 gate936 ( .A(N3137), .B(N2986), .Y(N3301) );
  OR2X1 gate937 ( .A(N3208), .B(N3029), .Y(N3302) );
  AND2X1 gate938 ( .A(N3172), .B(N3025), .Y(N3304) );
  AND2X1 gate939 ( .A(N3169), .B(N3022), .Y(N3306) );
  AND2X1 gate940 ( .A(N3166), .B(N3019), .Y(N3308) );
  AND2X1 gate941 ( .A(N3016), .B(N3163), .Y(N3309) );
  AND2X1 gate942 ( .A(N3160), .B(N3013), .Y(N3312) );
  AND2X1 gate943 ( .A(N3157), .B(N3010), .Y(N3314) );
  OR2X1 gate944 ( .A(N3215), .B(N3035), .Y(N3315) );
  OR2X1 gate945 ( .A(N3216), .B(N3036), .Y(N3318) );
  OR2X1 gate946 ( .A(N3217), .B(N3037), .Y(N3321) );
  OR2X1 gate947 ( .A(N3218), .B(N3044), .Y(N3324) );
  OR2X1 gate948 ( .A(N3219), .B(N3045), .Y(N3327) );
  OR2X1 gate949 ( .A(N3220), .B(N3046), .Y(N3330) );
  INVX1 gate950 ( .A(N3180), .Y(N3333) );
  OR2X1 gate951 ( .A(N3222), .B(N3053), .Y(N3334) );
  OR2X1 gate952 ( .A(N3223), .B(N3054), .Y(N3335) );
  OR2X1 gate953 ( .A(N3230), .B(N3064), .Y(N3336) );
  OR2X1 gate954 ( .A(N3231), .B(N3065), .Y(N3337) );
  BUFX2 gate955 ( .A(N3152), .Y(N3340) );
  BUFX2 gate956 ( .A(N3149), .Y(N3344) );
  BUFX2 gate957 ( .A(N3146), .Y(N3348) );
  BUFX2 gate958 ( .A(N3143), .Y(N3352) );
  BUFX2 gate959 ( .A(N3140), .Y(N3356) );
  BUFX2 gate960 ( .A(N3137), .Y(N3360) );
  BUFX2 gate961 ( .A(N3091), .Y(N3364) );
  BUFX2 gate962 ( .A(N3088), .Y(N3367) );
  BUFX2 gate963 ( .A(N3172), .Y(N3370) );
  BUFX2 gate964 ( .A(N3169), .Y(N3374) );
  BUFX2 gate965 ( .A(N3166), .Y(N3378) );
  BUFX2 gate966 ( .A(N3163), .Y(N3382) );
  BUFX2 gate967 ( .A(N3160), .Y(N3386) );
  BUFX2 gate968 ( .A(N3157), .Y(N3390) );
  BUFX2 gate969 ( .A(N3113), .Y(N3394) );
  BUFX2 gate970 ( .A(N3110), .Y(N3397) );
  NAND2X1 gate971 ( .A(N3195), .B(N3286), .Y(N3400) );
  NOR2X1 gate972 ( .A(N3281), .B(N3191), .Y(N3401) );
  NOR2X1 gate973 ( .A(N3282), .B(N3192), .Y(N3402) );
  NOR2X1 gate974 ( .A(N3283), .B(N3193), .Y(N3403) );
  NOR2X1 gate975 ( .A(N3284), .B(N3194), .Y(N3404) );
  INVX1 gate976 ( .A(N3238), .Y(N3405) );
  INVX1 gate977 ( .A(N3241), .Y(N3406) );
  AND2X1 gate978 ( .A(N3288), .B(N1836), .Y(N3409) );
  NAND2X1 gate979 ( .A(N2888), .B(N3333), .Y(N3410) );
  INVX1 gate980 ( .A(N3244), .Y(N3412) );
  INVX1 gate981 ( .A(N3247), .Y(N3414) );
  INVX1 gate982 ( .A(N3250), .Y(N3416) );
  INVX1 gate983 ( .A(N3253), .Y(N3418) );
  INVX1 gate984 ( .A(N3256), .Y(N3420) );
  INVX1 gate985 ( .A(N3259), .Y(N3422) );
  AND2X1 gate986 ( .A(N3302), .B(N1836), .Y(N3428) );
  INVX1 gate987 ( .A(N3262), .Y(N3430) );
  INVX1 gate988 ( .A(N3265), .Y(N3432) );
  INVX1 gate989 ( .A(N3268), .Y(N3434) );
  INVX1 gate990 ( .A(N3271), .Y(N3436) );
  INVX1 gate991 ( .A(N3274), .Y(N3438) );
  INVX1 gate992 ( .A(N3277), .Y(N3440) );
  AND2X1 gate993 ( .A(N3334), .B(N1190), .Y(N3450) );
  AND2X1 gate994 ( .A(N3335), .B(N1190), .Y(N3453) );
  AND2X1 gate995 ( .A(N3336), .B(N1195), .Y(N3456) );
  AND2X1 gate996 ( .A(N3337), .B(N1195), .Y(N3459) );
  AND2X1 gate997 ( .A(N3400), .B(N533), .Y(N3478) );
  AND2X1 gate998 ( .A(N3318), .B(N2128), .Y(N3479) );
  AND2X1 gate999 ( .A(N3315), .B(N1841), .Y(N3480) );
  NAND2X1 gate1000 ( .A(N3410), .B(N3289), .Y(N3481) );
  INVX1 gate1001 ( .A(N3340), .Y(N3482) );
  NAND2X1 gate1002 ( .A(N3340), .B(N3412), .Y(N3483) );
  INVX1 gate1003 ( .A(N3344), .Y(N3484) );
  NAND2X1 gate1004 ( .A(N3344), .B(N3414), .Y(N3485) );
  INVX1 gate1005 ( .A(N3348), .Y(N3486) );
  NAND2X1 gate1006 ( .A(N3348), .B(N3416), .Y(N3487) );
  INVX1 gate1007 ( .A(N3352), .Y(N3488) );
  NAND2X1 gate1008 ( .A(N3352), .B(N3418), .Y(N3489) );
  INVX1 gate1009 ( .A(N3356), .Y(N3490) );
  NAND2X1 gate1010 ( .A(N3356), .B(N3420), .Y(N3491) );
  INVX1 gate1011 ( .A(N3360), .Y(N3492) );
  NAND2X1 gate1012 ( .A(N3360), .B(N3422), .Y(N3493) );
  INVX1 gate1013 ( .A(N3364), .Y(N3494) );
  INVX1 gate1014 ( .A(N3367), .Y(N3496) );
  AND2X1 gate1015 ( .A(N3321), .B(N2135), .Y(N3498) );
  AND2X1 gate1016 ( .A(N3327), .B(N2128), .Y(N3499) );
  AND2X1 gate1017 ( .A(N3324), .B(N1841), .Y(N3500) );
  INVX1 gate1018 ( .A(N3370), .Y(N3501) );
  NAND2X1 gate1019 ( .A(N3370), .B(N3430), .Y(N3502) );
  INVX1 gate1020 ( .A(N3374), .Y(N3503) );
  NAND2X1 gate1021 ( .A(N3374), .B(N3432), .Y(N3504) );
  INVX1 gate1022 ( .A(N3378), .Y(N3505) );
  NAND2X1 gate1023 ( .A(N3378), .B(N3434), .Y(N3506) );
  INVX1 gate1024 ( .A(N3382), .Y(N3507) );
  NAND2X1 gate1025 ( .A(N3382), .B(N3436), .Y(N3508) );
  INVX1 gate1026 ( .A(N3386), .Y(N3509) );
  NAND2X1 gate1027 ( .A(N3386), .B(N3438), .Y(N3510) );
  INVX1 gate1028 ( .A(N3390), .Y(N3511) );
  NAND2X1 gate1029 ( .A(N3390), .B(N3440), .Y(N3512) );
  INVX1 gate1030 ( .A(N3394), .Y(N3513) );
  INVX1 gate1031 ( .A(N3397), .Y(N3515) );
  AND2X1 gate1032 ( .A(N3330), .B(N2135), .Y(N3517) );
  NAND2X1 gate1033 ( .A(N3402), .B(N3401), .Y(N3522) );
  NAND2X1 gate1034 ( .A(N3404), .B(N3403), .Y(N3525) );
  BUFX2 gate1035 ( .A(N3318), .Y(N3528) );
  BUFX2 gate1036 ( .A(N3315), .Y(N3531) );
  BUFX2 gate1037 ( .A(N3321), .Y(N3534) );
  BUFX2 gate1038 ( .A(N3327), .Y(N3537) );
  BUFX2 gate1039 ( .A(N3324), .Y(N3540) );
  BUFX2 gate1040 ( .A(N3330), .Y(N3543) );
  OR2X1 gate1041 ( .A(N3478), .B(N1813), .Y(N3546) );
  INVX1 gate1042 ( .A(N3481), .Y(N3551) );
  NAND2X1 gate1043 ( .A(N3244), .B(N3482), .Y(N3552) );
  NAND2X1 gate1044 ( .A(N3247), .B(N3484), .Y(N3553) );
  NAND2X1 gate1045 ( .A(N3250), .B(N3486), .Y(N3554) );
  NAND2X1 gate1046 ( .A(N3253), .B(N3488), .Y(N3555) );
  NAND2X1 gate1047 ( .A(N3256), .B(N3490), .Y(N3556) );
  NAND2X1 gate1048 ( .A(N3259), .B(N3492), .Y(N3557) );
  AND2X1 gate1049 ( .A(N3453), .B(N3091), .Y(N3558) );
  AND2X1 gate1050 ( .A(N3450), .B(N3088), .Y(N3559) );
  NAND2X1 gate1051 ( .A(N3262), .B(N3501), .Y(N3563) );
  NAND2X1 gate1052 ( .A(N3265), .B(N3503), .Y(N3564) );
  NAND2X1 gate1053 ( .A(N3268), .B(N3505), .Y(N3565) );
  NAND2X1 gate1054 ( .A(N3271), .B(N3507), .Y(N3566) );
  NAND2X1 gate1055 ( .A(N3274), .B(N3509), .Y(N3567) );
  NAND2X1 gate1056 ( .A(N3277), .B(N3511), .Y(N3568) );
  AND2X1 gate1057 ( .A(N3459), .B(N3113), .Y(N3569) );
  AND2X1 gate1058 ( .A(N3456), .B(N3110), .Y(N3570) );
  BUFX2 gate1059 ( .A(N3453), .Y(N3576) );
  BUFX2 gate1060 ( .A(N3450), .Y(N3579) );
  BUFX2 gate1061 ( .A(N3459), .Y(N3585) );
  BUFX2 gate1062 ( .A(N3456), .Y(N3588) );
  INVX1 gate1063 ( .A(N3522), .Y(N3592) );
  NAND2X1 gate1064 ( .A(N3522), .B(N3405), .Y(N3593) );
  INVX1 gate1065 ( .A(N3525), .Y(N3594) );
  NAND2X1 gate1066 ( .A(N3525), .B(N3406), .Y(N3595) );
  INVX1 gate1067 ( .A(N3528), .Y(N3596) );
  NAND2X1 gate1068 ( .A(N3528), .B(N2630), .Y(N3597) );
  NAND2X1 gate1069 ( .A(N3531), .B(N2376), .Y(N3598) );
  INVX1 gate1070 ( .A(N3531), .Y(N3599) );
  AND2X1 gate1071 ( .A(N3551), .B(N800), .Y(N3600) );
  NAND2X1 gate1072 ( .A(N3552), .B(N3483), .Y(N3603) );
  NAND2X1 gate1073 ( .A(N3553), .B(N3485), .Y(N3608) );
  NAND2X1 gate1074 ( .A(N3554), .B(N3487), .Y(N3612) );
  NAND2X1 gate1075 ( .A(N3555), .B(N3489), .Y(N3615) );
  NAND2X1 gate1076 ( .A(N3556), .B(N3491), .Y(N3616) );
  NAND2X1 gate1077 ( .A(N3557), .B(N3493), .Y(N3622) );
  INVX1 gate1078 ( .A(N3534), .Y(N3629) );
  NAND2X1 gate1079 ( .A(N3534), .B(N2645), .Y(N3630) );
  INVX1 gate1080 ( .A(N3537), .Y(N3631) );
  NAND2X1 gate1081 ( .A(N3537), .B(N2655), .Y(N3632) );
  NAND2X1 gate1082 ( .A(N3540), .B(N2403), .Y(N3633) );
  INVX1 gate1083 ( .A(N3540), .Y(N3634) );
  NAND2X1 gate1084 ( .A(N3563), .B(N3502), .Y(N3635) );
  NAND2X1 gate1085 ( .A(N3564), .B(N3504), .Y(N3640) );
  NAND2X1 gate1086 ( .A(N3565), .B(N3506), .Y(N3644) );
  NAND2X1 gate1087 ( .A(N3566), .B(N3508), .Y(N3647) );
  NAND2X1 gate1088 ( .A(N3567), .B(N3510), .Y(N3648) );
  NAND2X1 gate1089 ( .A(N3568), .B(N3512), .Y(N3654) );
  INVX1 gate1090 ( .A(N3543), .Y(N3661) );
  NAND2X1 gate1091 ( .A(N3543), .B(N2656), .Y(N3662) );
  NAND2X1 gate1092 ( .A(N3238), .B(N3592), .Y(N3667) );
  NAND2X1 gate1093 ( .A(N3241), .B(N3594), .Y(N3668) );
  NAND2X1 gate1094 ( .A(N2472), .B(N3596), .Y(N3669) );
  NAND2X1 gate1095 ( .A(N2213), .B(N3599), .Y(N3670) );
  BUFX2 gate1096 ( .A(N3600), .Y(N3671) );
  INVX1 gate1097 ( .A(N3576), .Y(N3691) );
  NAND2X1 gate1098 ( .A(N3576), .B(N3494), .Y(N3692) );
  INVX1 gate1099 ( .A(N3579), .Y(N3693) );
  NAND2X1 gate1100 ( .A(N3579), .B(N3496), .Y(N3694) );
  NAND2X1 gate1101 ( .A(N2475), .B(N3629), .Y(N3695) );
  NAND2X1 gate1102 ( .A(N2478), .B(N3631), .Y(N3696) );
  NAND2X1 gate1103 ( .A(N2216), .B(N3634), .Y(N3697) );
  INVX1 gate1104 ( .A(N3585), .Y(N3716) );
  NAND2X1 gate1105 ( .A(N3585), .B(N3513), .Y(N3717) );
  INVX1 gate1106 ( .A(N3588), .Y(N3718) );
  NAND2X1 gate1107 ( .A(N3588), .B(N3515), .Y(N3719) );
  NAND2X1 gate1108 ( .A(N2481), .B(N3661), .Y(N3720) );
  NAND2X1 gate1109 ( .A(N3667), .B(N3593), .Y(N3721) );
  NAND2X1 gate1110 ( .A(N3668), .B(N3595), .Y(N3722) );
  NAND2X1 gate1111 ( .A(N3669), .B(N3597), .Y(N3723) );
  NAND2X1 gate1112 ( .A(N3670), .B(N3598), .Y(N3726) );
  INVX1 gate1113 ( .A(N3600), .Y(N3727) );
  NAND2X1 gate1114 ( .A(N3364), .B(N3691), .Y(N3728) );
  NAND2X1 gate1115 ( .A(N3367), .B(N3693), .Y(N3729) );
  NAND2X1 gate1116 ( .A(N3695), .B(N3630), .Y(N3730) );
  AND2X1 gate1117_1 ( .A(N3608), .B(N3615), .Y(N3731_1) );
  AND2X1 gate1117_2 ( .A(N3612), .B(N3603), .Y(N3731_2) );
  AND2X1 gate1117 ( .A(N3731_1), .B(N3731_2), .Y(N3731) );
  AND2X1 gate1118 ( .A(N3603), .B(N3293), .Y(N3732) );
  AND2X1 gate1119_1 ( .A(N3608), .B(N3603), .Y(N3733_1) );
  AND2X1 gate1119 ( .A(N3295), .B(N3733_1), .Y(N3733) );
  AND2X1 gate1120_1 ( .A(N3612), .B(N3603), .Y(N3734_1) );
  AND2X1 gate1120_2 ( .A(N3296), .B(N3608), .Y(N3734_2) );
  AND2X1 gate1120 ( .A(N3734_1), .B(N3734_2), .Y(N3734) );
  AND2X1 gate1121 ( .A(N3616), .B(N3301), .Y(N3735) );
  AND2X1 gate1122_1 ( .A(N3622), .B(N3616), .Y(N3736_1) );
  AND2X1 gate1122 ( .A(N3558), .B(N3736_1), .Y(N3736) );
  NAND2X1 gate1123 ( .A(N3696), .B(N3632), .Y(N3737) );
  NAND2X1 gate1124 ( .A(N3697), .B(N3633), .Y(N3740) );
  NAND2X1 gate1125 ( .A(N3394), .B(N3716), .Y(N3741) );
  NAND2X1 gate1126 ( .A(N3397), .B(N3718), .Y(N3742) );
  NAND2X1 gate1127 ( .A(N3720), .B(N3662), .Y(N3743) );
  AND2X1 gate1128_1 ( .A(N3640), .B(N3647), .Y(N3744_1) );
  AND2X1 gate1128_2 ( .A(N3644), .B(N3635), .Y(N3744_2) );
  AND2X1 gate1128 ( .A(N3744_1), .B(N3744_2), .Y(N3744) );
  AND2X1 gate1129 ( .A(N3635), .B(N3306), .Y(N3745) );
  AND2X1 gate1130_1 ( .A(N3640), .B(N3635), .Y(N3746_1) );
  AND2X1 gate1130 ( .A(N3308), .B(N3746_1), .Y(N3746) );
  AND2X1 gate1131_1 ( .A(N3644), .B(N3635), .Y(N3747_1) );
  AND2X1 gate1131_2 ( .A(N3309), .B(N3640), .Y(N3747_2) );
  AND2X1 gate1131 ( .A(N3747_1), .B(N3747_2), .Y(N3747) );
  AND2X1 gate1132 ( .A(N3648), .B(N3314), .Y(N3748) );
  AND2X1 gate1133_1 ( .A(N3654), .B(N3648), .Y(N3749_1) );
  AND2X1 gate1133 ( .A(N3569), .B(N3749_1), .Y(N3749) );
  INVX1 gate1134 ( .A(N3721), .Y(N3750) );
  AND2X1 gate1135 ( .A(N3722), .B(N246), .Y(N3753) );
  NAND2X1 gate1136 ( .A(N3728), .B(N3692), .Y(N3754) );
  NAND2X1 gate1137 ( .A(N3729), .B(N3694), .Y(N3758) );
  INVX1 gate1138 ( .A(N3731), .Y(N3761) );
  OR2X1 gate1139_1 ( .A(N3291), .B(N3732), .Y(N3762_1) );
  OR2X1 gate1139_2 ( .A(N3733), .B(N3734), .Y(N3762_2) );
  OR2X1 gate1139 ( .A(N3762_1), .B(N3762_2), .Y(N3762) );
  NAND2X1 gate1140 ( .A(N3741), .B(N3717), .Y(N3767) );
  NAND2X1 gate1141 ( .A(N3742), .B(N3719), .Y(N3771) );
  INVX1 gate1142 ( .A(N3744), .Y(N3774) );
  OR2X1 gate1143_1 ( .A(N3304), .B(N3745), .Y(N3775_1) );
  OR2X1 gate1143_2 ( .A(N3746), .B(N3747), .Y(N3775_2) );
  OR2X1 gate1143 ( .A(N3775_1), .B(N3775_2), .Y(N3775) );
  AND2X1 gate1144 ( .A(N3723), .B(N3480), .Y(N3778) );
  AND2X1 gate1145_1 ( .A(N3726), .B(N3723), .Y(N3779_1) );
  AND2X1 gate1145 ( .A(N3409), .B(N3779_1), .Y(N3779) );
  OR2X1 gate1146 ( .A(N2125), .B(N3753), .Y(N3780) );
  AND2X1 gate1147 ( .A(N3750), .B(N800), .Y(N3790) );
  AND2X1 gate1148 ( .A(N3737), .B(N3500), .Y(N3793) );
  AND2X1 gate1149_1 ( .A(N3740), .B(N3737), .Y(N3794_1) );
  AND2X1 gate1149 ( .A(N3428), .B(N3794_1), .Y(N3794) );
  OR2X1 gate1150_1 ( .A(N3479), .B(N3778), .Y(N3802_1) );
  OR2X1 gate1150 ( .A(N3779), .B(N3802_1), .Y(N3802) );
  BUFX2 gate1151 ( .A(N3780), .Y(N3803) );
  BUFX2 gate1152 ( .A(N3780), .Y(N3804) );
  INVX1 gate1153 ( .A(N3762), .Y(N3805) );
  AND2X1 gate1154_1 ( .A(N3622), .B(N3730), .Y(N3806_1) );
  AND2X1 gate1154_2 ( .A(N3754), .B(N3616), .Y(N3806_2) );
  AND2X1 gate1154_3 ( .A(N3758), .B(N3806_1), .Y(N3806_3) );
  AND2X1 gate1154 ( .A(N3806_2), .B(N3806_3), .Y(N3806) );
  AND2X1 gate1155_1 ( .A(N3754), .B(N3616), .Y(N3807_1) );
  AND2X1 gate1155_2 ( .A(N3559), .B(N3622), .Y(N3807_2) );
  AND2X1 gate1155 ( .A(N3807_1), .B(N3807_2), .Y(N3807) );
  AND2X1 gate1156_1 ( .A(N3758), .B(N3754), .Y(N3808_1) );
  AND2X1 gate1156_2 ( .A(N3616), .B(N3498), .Y(N3808_2) );
  AND2X1 gate1156_3 ( .A(N3622), .B(N3808_1), .Y(N3808_3) );
  AND2X1 gate1156 ( .A(N3808_2), .B(N3808_3), .Y(N3808) );
  BUFX2 gate1157 ( .A(N3790), .Y(N3809) );
  OR2X1 gate1158_1 ( .A(N3499), .B(N3793), .Y(N3811_1) );
  OR2X1 gate1158 ( .A(N3794), .B(N3811_1), .Y(N3811) );
  INVX1 gate1159 ( .A(N3775), .Y(N3812) );
  AND2X1 gate1160_1 ( .A(N3654), .B(N3743), .Y(N3813_1) );
  AND2X1 gate1160_2 ( .A(N3767), .B(N3648), .Y(N3813_2) );
  AND2X1 gate1160_3 ( .A(N3771), .B(N3813_1), .Y(N3813_3) );
  AND2X1 gate1160 ( .A(N3813_2), .B(N3813_3), .Y(N3813) );
  AND2X1 gate1161_1 ( .A(N3767), .B(N3648), .Y(N3814_1) );
  AND2X1 gate1161_2 ( .A(N3570), .B(N3654), .Y(N3814_2) );
  AND2X1 gate1161 ( .A(N3814_1), .B(N3814_2), .Y(N3814) );
  AND2X1 gate1162_1 ( .A(N3771), .B(N3767), .Y(N3815_1) );
  AND2X1 gate1162_2 ( .A(N3648), .B(N3517), .Y(N3815_2) );
  AND2X1 gate1162_3 ( .A(N3654), .B(N3815_1), .Y(N3815_3) );
  AND2X1 gate1162 ( .A(N3815_2), .B(N3815_3), .Y(N3815) );
  OR2X1 gate1163_1 ( .A(N3299), .B(N3735), .Y(N3816_1) );
  OR2X1 gate1163_2 ( .A(N3736), .B(N3807), .Y(N3816_2) );
  OR2X1 gate1163_3 ( .A(N3808), .B(N3816_1), .Y(N3816_3) );
  OR2X1 gate1163 ( .A(N3816_2), .B(N3816_3), .Y(N3816) );
  AND2X1 gate1164 ( .A(N3806), .B(N3802), .Y(N3817) );
  NAND2X1 gate1165 ( .A(N3805), .B(N3761), .Y(N3818) );
  INVX1 gate1166 ( .A(N3790), .Y(N3819) );
  OR2X1 gate1167_1 ( .A(N3312), .B(N3748), .Y(N3820_1) );
  OR2X1 gate1167_2 ( .A(N3749), .B(N3814), .Y(N3820_2) );
  OR2X1 gate1167_3 ( .A(N3815), .B(N3820_1), .Y(N3820_3) );
  OR2X1 gate1167 ( .A(N3820_2), .B(N3820_3), .Y(N3820) );
  AND2X1 gate1168 ( .A(N3813), .B(N3811), .Y(N3821) );
  NAND2X1 gate1169 ( .A(N3812), .B(N3774), .Y(N3822) );
  OR2X1 gate1170 ( .A(N3816), .B(N3817), .Y(N3823) );
  AND2X1 gate1171_1 ( .A(N3727), .B(N3819), .Y(N3826_1) );
  AND2X1 gate1171 ( .A(N2841), .B(N3826_1), .Y(N3826) );
  OR2X1 gate1172 ( .A(N3820), .B(N3821), .Y(N3827) );
  INVX1 gate1173 ( .A(N3823), .Y(N3834) );
  AND2X1 gate1174 ( .A(N3818), .B(N3823), .Y(N3835) );
  INVX1 gate1175 ( .A(N3827), .Y(N3836) );
  AND2X1 gate1176 ( .A(N3822), .B(N3827), .Y(N3837) );
  AND2X1 gate1177 ( .A(N3762), .B(N3834), .Y(N3838) );
  AND2X1 gate1178 ( .A(N3775), .B(N3836), .Y(N3839) );
  OR2X1 gate1179 ( .A(N3838), .B(N3835), .Y(N3840) );
  OR2X1 gate1180 ( .A(N3839), .B(N3837), .Y(N3843) );
  BUFX2 gate1181 ( .A(N3843), .Y(N3851) );
  NAND2X1 gate1182 ( .A(N3843), .B(N3840), .Y(N3852) );
  AND2X1 gate1183 ( .A(N3843), .B(N3852), .Y(N3857) );
  AND2X1 gate1184 ( .A(N3852), .B(N3840), .Y(N3858) );
  OR2X1 gate1185 ( .A(N3857), .B(N3858), .Y(N3859) );
  INVX1 gate1186 ( .A(N3859), .Y(N3864) );
  AND2X1 gate1187 ( .A(N3859), .B(N3864), .Y(N3869) );
  OR2X1 gate1188 ( .A(N3869), .B(N3864), .Y(N3870) );
  INVX1 gate1189 ( .A(N3870), .Y(N3875) );
  AND2X1 gate1190_1 ( .A(N2826), .B(N3028), .Y(N3876_1) );
  AND2X1 gate1190 ( .A(N3870), .B(N3876_1), .Y(N3876) );
  AND2X1 gate1191_1 ( .A(N3826), .B(N3876), .Y(N3877_1) );
  AND2X1 gate1191 ( .A(N1591), .B(N3877_1), .Y(N3877) );
  BUFX2 gate1192 ( .A(N3877), .Y(N3881) );
  INVX1 gate1193 ( .A(N3877), .Y(N3882) );
  BUFX2 gate1194 ( .A(N143_I), .Y(N143_O) );
  BUFX2 gate1195 ( .A(N144_I), .Y(N144_O) );
  BUFX2 gate1196 ( .A(N145_I), .Y(N145_O) );
  BUFX2 gate1197 ( .A(N146_I), .Y(N146_O) );
  BUFX2 gate1198 ( .A(N147_I), .Y(N147_O) );
  BUFX2 gate1199 ( .A(N148_I), .Y(N148_O) );
  BUFX2 gate1200 ( .A(N149_I), .Y(N149_O) );
  BUFX2 gate1201 ( .A(N150_I), .Y(N150_O) );
  BUFX2 gate1202 ( .A(N151_I), .Y(N151_O) );
  BUFX2 gate1203 ( .A(N152_I), .Y(N152_O) );
  BUFX2 gate1204 ( .A(N153_I), .Y(N153_O) );
  BUFX2 gate1205 ( .A(N154_I), .Y(N154_O) );
  BUFX2 gate1206 ( .A(N155_I), .Y(N155_O) );
  BUFX2 gate1207 ( .A(N156_I), .Y(N156_O) );
  BUFX2 gate1208 ( .A(N157_I), .Y(N157_O) );
  BUFX2 gate1209 ( .A(N158_I), .Y(N158_O) );
  BUFX2 gate1210 ( .A(N159_I), .Y(N159_O) );
  BUFX2 gate1211 ( .A(N160_I), .Y(N160_O) );
  BUFX2 gate1212 ( .A(N161_I), .Y(N161_O) );
  BUFX2 gate1213 ( .A(N162_I), .Y(N162_O) );
  BUFX2 gate1214 ( .A(N163_I), .Y(N163_O) );
  BUFX2 gate1215 ( .A(N164_I), .Y(N164_O) );
  BUFX2 gate1216 ( .A(N165_I), .Y(N165_O) );
  BUFX2 gate1217 ( .A(N166_I), .Y(N166_O) );
  BUFX2 gate1218 ( .A(N167_I), .Y(N167_O) );
  BUFX2 gate1219 ( .A(N168_I), .Y(N168_O) );
  BUFX2 gate1220 ( .A(N169_I), .Y(N169_O) );
  BUFX2 gate1221 ( .A(N170_I), .Y(N170_O) );
  BUFX2 gate1222 ( .A(N171_I), .Y(N171_O) );
  BUFX2 gate1223 ( .A(N172_I), .Y(N172_O) );
  BUFX2 gate1224 ( .A(N173_I), .Y(N173_O) );
  BUFX2 gate1225 ( .A(N174_I), .Y(N174_O) );
  BUFX2 gate1226 ( .A(N175_I), .Y(N175_O) );
  BUFX2 gate1227 ( .A(N176_I), .Y(N176_O) );
  BUFX2 gate1228 ( .A(N177_I), .Y(N177_O) );
  BUFX2 gate1229 ( .A(N178_I), .Y(N178_O) );
  BUFX2 gate1230 ( .A(N179_I), .Y(N179_O) );
  BUFX2 gate1231 ( .A(N180_I), .Y(N180_O) );
  BUFX2 gate1232 ( .A(N181_I), .Y(N181_O) );
  BUFX2 gate1233 ( .A(N182_I), .Y(N182_O) );
  BUFX2 gate1234 ( .A(N183_I), .Y(N183_O) );
  BUFX2 gate1235 ( .A(N184_I), .Y(N184_O) );
  BUFX2 gate1236 ( .A(N185_I), .Y(N185_O) );
  BUFX2 gate1237 ( .A(N186_I), .Y(N186_O) );
  BUFX2 gate1238 ( .A(N187_I), .Y(N187_O) );
  BUFX2 gate1239 ( .A(N188_I), .Y(N188_O) );
  BUFX2 gate1240 ( .A(N189_I), .Y(N189_O) );
  BUFX2 gate1241 ( .A(N190_I), .Y(N190_O) );
  BUFX2 gate1242 ( .A(N191_I), .Y(N191_O) );
  BUFX2 gate1243 ( .A(N192_I), .Y(N192_O) );
  BUFX2 gate1244 ( .A(N193_I), .Y(N193_O) );
  BUFX2 gate1245 ( .A(N194_I), .Y(N194_O) );
  BUFX2 gate1246 ( .A(N195_I), .Y(N195_O) );
  BUFX2 gate1247 ( .A(N196_I), .Y(N196_O) );
  BUFX2 gate1248 ( .A(N197_I), .Y(N197_O) );
  BUFX2 gate1249 ( .A(N198_I), .Y(N198_O) );
  BUFX2 gate1250 ( .A(N199_I), .Y(N199_O) );
  BUFX2 gate1251 ( .A(N200_I), .Y(N200_O) );
  BUFX2 gate1252 ( .A(N201_I), .Y(N201_O) );
  BUFX2 gate1253 ( .A(N202_I), .Y(N202_O) );
  BUFX2 gate1254 ( .A(N203_I), .Y(N203_O) );
  BUFX2 gate1255 ( .A(N204_I), .Y(N204_O) );
  BUFX2 gate1256 ( .A(N205_I), .Y(N205_O) );
  BUFX2 gate1257 ( .A(N206_I), .Y(N206_O) );
  BUFX2 gate1258 ( .A(N207_I), .Y(N207_O) );
  BUFX2 gate1259 ( .A(N208_I), .Y(N208_O) );
  BUFX2 gate1260 ( .A(N209_I), .Y(N209_O) );
  BUFX2 gate1261 ( .A(N210_I), .Y(N210_O) );
  BUFX2 gate1262 ( .A(N211_I), .Y(N211_O) );
  BUFX2 gate1263 ( .A(N212_I), .Y(N212_O) );
  BUFX2 gate1264 ( .A(N213_I), .Y(N213_O) );
  BUFX2 gate1265 ( .A(N214_I), .Y(N214_O) );
  BUFX2 gate1266 ( .A(N215_I), .Y(N215_O) );
  BUFX2 gate1267 ( .A(N216_I), .Y(N216_O) );
  BUFX2 gate1268 ( .A(N217_I), .Y(N217_O) );
  BUFX2 gate1269 ( .A(N218_I), .Y(N218_O) );
endmodule

